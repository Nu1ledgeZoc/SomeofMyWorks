module rom3 (
    clk,
    otp
);
    input clk;
    output reg[7:0]otp;
    reg [7:0] data[999:0];
    reg [9:0] count;
    reg [9:0] mod;
    initial begin
         count=0;
        mod=1000;
        data[999]=0;
        data[998]=1;
        data[997]=1;
        data[996]=2;
        data[995]=2;
        data[994]=3;
        data[993]=3;
        data[992]=4;
        data[991]=4;
        data[990]=5;
        data[989]=5;
        data[988]=6;
        data[987]=6;
        data[986]=7;
        data[985]=7;
        data[984]=8;
        data[983]=8;
        data[982]=9;
        data[981]=9;
        data[980]=10;
        data[979]=10;
        data[978]=11;
        data[977]=11;
        data[976]=12;
        data[975]=12;
        data[974]=13;
        data[973]=13;
        data[972]=14;
        data[971]=14;
        data[970]=15;
        data[969]=15;
        data[968]=16;
        data[967]=16;
        data[966]=17;
        data[965]=17;
        data[964]=18;
        data[963]=18;
        data[962]=19;
        data[961]=19;
        data[960]=20;
        data[959]=20;
        data[958]=21;
        data[957]=21;
        data[956]=22;
        data[955]=22;
        data[954]=23;
        data[953]=23;
        data[952]=24;
        data[951]=24;
        data[950]=25;
        data[949]=25;
        data[948]=26;
        data[947]=27;
        data[946]=27;
        data[945]=28;
        data[944]=28;
        data[943]=29;
        data[942]=29;
        data[941]=30;
        data[940]=30;
        data[939]=31;
        data[938]=31;
        data[937]=32;
        data[936]=32;
        data[935]=33;
        data[934]=33;
        data[933]=34;
        data[932]=34;
        data[931]=35;
        data[930]=35;
        data[929]=36;
        data[928]=36;
        data[927]=37;
        data[926]=37;
        data[925]=38;
        data[924]=38;
        data[923]=39;
        data[922]=39;
        data[921]=40;
        data[920]=40;
        data[919]=41;
        data[918]=41;
        data[917]=42;
        data[916]=42;
        data[915]=43;
        data[914]=43;
        data[913]=44;
        data[912]=44;
        data[911]=45;
        data[910]=45;
        data[909]=46;
        data[908]=46;
        data[907]=47;
        data[906]=47;
        data[905]=48;
        data[904]=48;
        data[903]=49;
        data[902]=49;
        data[901]=50;
        data[900]=50;
        data[899]=51;
        data[898]=52;
        data[897]=52;
        data[896]=53;
        data[895]=53;
        data[894]=54;
        data[893]=54;
        data[892]=55;
        data[891]=55;
        data[890]=56;
        data[889]=56;
        data[888]=57;
        data[887]=57;
        data[886]=58;
        data[885]=58;
        data[884]=59;
        data[883]=59;
        data[882]=60;
        data[881]=60;
        data[880]=61;
        data[879]=61;
        data[878]=62;
        data[877]=62;
        data[876]=63;
        data[875]=63;
        data[874]=64;
        data[873]=64;
        data[872]=65;
        data[871]=65;
        data[870]=66;
        data[869]=66;
        data[868]=67;
        data[867]=67;
        data[866]=68;
        data[865]=68;
        data[864]=69;
        data[863]=69;
        data[862]=70;
        data[861]=70;
        data[860]=71;
        data[859]=71;
        data[858]=72;
        data[857]=72;
        data[856]=73;
        data[855]=73;
        data[854]=74;
        data[853]=74;
        data[852]=75;
        data[851]=75;
        data[850]=76;
        data[849]=77;
        data[848]=77;
        data[847]=78;
        data[846]=78;
        data[845]=79;
        data[844]=79;
        data[843]=80;
        data[842]=80;
        data[841]=81;
        data[840]=81;
        data[839]=82;
        data[838]=82;
        data[837]=83;
        data[836]=83;
        data[835]=84;
        data[834]=84;
        data[833]=85;
        data[832]=85;
        data[831]=86;
        data[830]=86;
        data[829]=87;
        data[828]=87;
        data[827]=88;
        data[826]=88;
        data[825]=89;
        data[824]=89;
        data[823]=90;
        data[822]=90;
        data[821]=91;
        data[820]=91;
        data[819]=92;
        data[818]=92;
        data[817]=93;
        data[816]=93;
        data[815]=94;
        data[814]=94;
        data[813]=95;
        data[812]=95;
        data[811]=96;
        data[810]=96;
        data[809]=97;
        data[808]=97;
        data[807]=98;
        data[806]=98;
        data[805]=99;
        data[804]=99;
        data[803]=100;
        data[802]=100;
        data[801]=101;
        data[800]=101;
        data[799]=102;
        data[798]=103;
        data[797]=103;
        data[796]=104;
        data[795]=104;
        data[794]=105;
        data[793]=105;
        data[792]=106;
        data[791]=106;
        data[790]=107;
        data[789]=107;
        data[788]=108;
        data[787]=108;
        data[786]=109;
        data[785]=109;
        data[784]=110;
        data[783]=110;
        data[782]=111;
        data[781]=111;
        data[780]=112;
        data[779]=112;
        data[778]=113;
        data[777]=113;
        data[776]=114;
        data[775]=114;
        data[774]=115;
        data[773]=115;
        data[772]=116;
        data[771]=116;
        data[770]=117;
        data[769]=117;
        data[768]=118;
        data[767]=118;
        data[766]=119;
        data[765]=119;
        data[764]=120;
        data[763]=120;
        data[762]=121;
        data[761]=121;
        data[760]=122;
        data[759]=122;
        data[758]=123;
        data[757]=123;
        data[756]=124;
        data[755]=124;
        data[754]=125;
        data[753]=125;
        data[752]=126;
        data[751]=126;
        data[750]=127;
        data[749]=128;
        data[748]=128;
        data[747]=129;
        data[746]=129;
        data[745]=130;
        data[744]=130;
        data[743]=131;
        data[742]=131;
        data[741]=132;
        data[740]=132;
        data[739]=133;
        data[738]=133;
        data[737]=134;
        data[736]=134;
        data[735]=135;
        data[734]=135;
        data[733]=136;
        data[732]=136;
        data[731]=137;
        data[730]=137;
        data[729]=138;
        data[728]=138;
        data[727]=139;
        data[726]=139;
        data[725]=140;
        data[724]=140;
        data[723]=141;
        data[722]=141;
        data[721]=142;
        data[720]=142;
        data[719]=143;
        data[718]=143;
        data[717]=144;
        data[716]=144;
        data[715]=145;
        data[714]=145;
        data[713]=146;
        data[712]=146;
        data[711]=147;
        data[710]=147;
        data[709]=148;
        data[708]=148;
        data[707]=149;
        data[706]=149;
        data[705]=150;
        data[704]=150;
        data[703]=151;
        data[702]=151;
        data[701]=152;
        data[700]=152;
        data[699]=153;
        data[698]=154;
        data[697]=154;
        data[696]=155;
        data[695]=155;
        data[694]=156;
        data[693]=156;
        data[692]=157;
        data[691]=157;
        data[690]=158;
        data[689]=158;
        data[688]=159;
        data[687]=159;
        data[686]=160;
        data[685]=160;
        data[684]=161;
        data[683]=161;
        data[682]=162;
        data[681]=162;
        data[680]=163;
        data[679]=163;
        data[678]=164;
        data[677]=164;
        data[676]=165;
        data[675]=165;
        data[674]=166;
        data[673]=166;
        data[672]=167;
        data[671]=167;
        data[670]=168;
        data[669]=168;
        data[668]=169;
        data[667]=169;
        data[666]=170;
        data[665]=170;
        data[664]=171;
        data[663]=171;
        data[662]=172;
        data[661]=172;
        data[660]=173;
        data[659]=173;
        data[658]=174;
        data[657]=174;
        data[656]=175;
        data[655]=175;
        data[654]=176;
        data[653]=176;
        data[652]=177;
        data[651]=177;
        data[650]=178;
        data[649]=179;
        data[648]=179;
        data[647]=180;
        data[646]=180;
        data[645]=181;
        data[644]=181;
        data[643]=182;
        data[642]=182;
        data[641]=183;
        data[640]=183;
        data[639]=184;
        data[638]=184;
        data[637]=185;
        data[636]=185;
        data[635]=186;
        data[634]=186;
        data[633]=187;
        data[632]=187;
        data[631]=188;
        data[630]=188;
        data[629]=189;
        data[628]=189;
        data[627]=190;
        data[626]=190;
        data[625]=191;
        data[624]=191;
        data[623]=192;
        data[622]=192;
        data[621]=193;
        data[620]=193;
        data[619]=194;
        data[618]=194;
        data[617]=195;
        data[616]=195;
        data[615]=196;
        data[614]=196;
        data[613]=197;
        data[612]=197;
        data[611]=198;
        data[610]=198;
        data[609]=199;
        data[608]=199;
        data[607]=200;
        data[606]=200;
        data[605]=201;
        data[604]=201;
        data[603]=202;
        data[602]=202;
        data[601]=203;
        data[600]=203;
        data[599]=204;
        data[598]=205;
        data[597]=205;
        data[596]=206;
        data[595]=206;
        data[594]=207;
        data[593]=207;
        data[592]=208;
        data[591]=208;
        data[590]=209;
        data[589]=209;
        data[588]=210;
        data[587]=210;
        data[586]=211;
        data[585]=211;
        data[584]=212;
        data[583]=212;
        data[582]=213;
        data[581]=213;
        data[580]=214;
        data[579]=214;
        data[578]=215;
        data[577]=215;
        data[576]=216;
        data[575]=216;
        data[574]=217;
        data[573]=217;
        data[572]=218;
        data[571]=218;
        data[570]=219;
        data[569]=219;
        data[568]=220;
        data[567]=220;
        data[566]=221;
        data[565]=221;
        data[564]=222;
        data[563]=222;
        data[562]=223;
        data[561]=223;
        data[560]=224;
        data[559]=224;
        data[558]=225;
        data[557]=225;
        data[556]=226;
        data[555]=226;
        data[554]=227;
        data[553]=227;
        data[552]=228;
        data[551]=228;
        data[550]=229;
        data[549]=230;
        data[548]=230;
        data[547]=231;
        data[546]=231;
        data[545]=232;
        data[544]=232;
        data[543]=233;
        data[542]=233;
        data[541]=234;
        data[540]=234;
        data[539]=235;
        data[538]=235;
        data[537]=236;
        data[536]=236;
        data[535]=237;
        data[534]=237;
        data[533]=238;
        data[532]=238;
        data[531]=239;
        data[530]=239;
        data[529]=240;
        data[528]=240;
        data[527]=241;
        data[526]=241;
        data[525]=242;
        data[524]=242;
        data[523]=243;
        data[522]=243;
        data[521]=244;
        data[520]=244;
        data[519]=245;
        data[518]=245;
        data[517]=246;
        data[516]=246;
        data[515]=247;
        data[514]=247;
        data[513]=248;
        data[512]=248;
        data[511]=249;
        data[510]=249;
        data[509]=250;
        data[508]=250;
        data[507]=251;
        data[506]=251;
        data[505]=252;
        data[504]=252;
        data[503]=253;
        data[502]=253;
        data[501]=254;
        data[500]=254;
        data[499]=254;
        data[498]=254;
        data[497]=253;
        data[496]=253;
        data[495]=252;
        data[494]=252;
        data[493]=251;
        data[492]=251;
        data[491]=250;
        data[490]=250;
        data[489]=249;
        data[488]=249;
        data[487]=248;
        data[486]=248;
        data[485]=247;
        data[484]=247;
        data[483]=246;
        data[482]=246;
        data[481]=245;
        data[480]=245;
        data[479]=244;
        data[478]=244;
        data[477]=243;
        data[476]=243;
        data[475]=242;
        data[474]=242;
        data[473]=241;
        data[472]=241;
        data[471]=240;
        data[470]=240;
        data[469]=239;
        data[468]=239;
        data[467]=238;
        data[466]=238;
        data[465]=237;
        data[464]=237;
        data[463]=236;
        data[462]=236;
        data[461]=235;
        data[460]=235;
        data[459]=234;
        data[458]=234;
        data[457]=233;
        data[456]=233;
        data[455]=232;
        data[454]=232;
        data[453]=231;
        data[452]=231;
        data[451]=230;
        data[450]=230;
        data[449]=229;
        data[448]=228;
        data[447]=228;
        data[446]=227;
        data[445]=227;
        data[444]=226;
        data[443]=226;
        data[442]=225;
        data[441]=225;
        data[440]=224;
        data[439]=224;
        data[438]=223;
        data[437]=223;
        data[436]=222;
        data[435]=222;
        data[434]=221;
        data[433]=221;
        data[432]=220;
        data[431]=220;
        data[430]=219;
        data[429]=219;
        data[428]=218;
        data[427]=218;
        data[426]=217;
        data[425]=217;
        data[424]=216;
        data[423]=216;
        data[422]=215;
        data[421]=215;
        data[420]=214;
        data[419]=214;
        data[418]=213;
        data[417]=213;
        data[416]=212;
        data[415]=212;
        data[414]=211;
        data[413]=211;
        data[412]=210;
        data[411]=210;
        data[410]=209;
        data[409]=209;
        data[408]=208;
        data[407]=208;
        data[406]=207;
        data[405]=207;
        data[404]=206;
        data[403]=206;
        data[402]=205;
        data[401]=205;
        data[400]=204;
        data[399]=203;
        data[398]=203;
        data[397]=202;
        data[396]=202;
        data[395]=201;
        data[394]=201;
        data[393]=200;
        data[392]=200;
        data[391]=199;
        data[390]=199;
        data[389]=198;
        data[388]=198;
        data[387]=197;
        data[386]=197;
        data[385]=196;
        data[384]=196;
        data[383]=195;
        data[382]=195;
        data[381]=194;
        data[380]=194;
        data[379]=193;
        data[378]=193;
        data[377]=192;
        data[376]=192;
        data[375]=191;
        data[374]=191;
        data[373]=190;
        data[372]=190;
        data[371]=189;
        data[370]=189;
        data[369]=188;
        data[368]=188;
        data[367]=187;
        data[366]=187;
        data[365]=186;
        data[364]=186;
        data[363]=185;
        data[362]=185;
        data[361]=184;
        data[360]=184;
        data[359]=183;
        data[358]=183;
        data[357]=182;
        data[356]=182;
        data[355]=181;
        data[354]=181;
        data[353]=180;
        data[352]=180;
        data[351]=179;
        data[350]=179;
        data[349]=178;
        data[348]=177;
        data[347]=177;
        data[346]=176;
        data[345]=176;
        data[344]=175;
        data[343]=175;
        data[342]=174;
        data[341]=174;
        data[340]=173;
        data[339]=173;
        data[338]=172;
        data[337]=172;
        data[336]=171;
        data[335]=171;
        data[334]=170;
        data[333]=170;
        data[332]=169;
        data[331]=169;
        data[330]=168;
        data[329]=168;
        data[328]=167;
        data[327]=167;
        data[326]=166;
        data[325]=166;
        data[324]=165;
        data[323]=165;
        data[322]=164;
        data[321]=164;
        data[320]=163;
        data[319]=163;
        data[318]=162;
        data[317]=162;
        data[316]=161;
        data[315]=161;
        data[314]=160;
        data[313]=160;
        data[312]=159;
        data[311]=159;
        data[310]=158;
        data[309]=158;
        data[308]=157;
        data[307]=157;
        data[306]=156;
        data[305]=156;
        data[304]=155;
        data[303]=155;
        data[302]=154;
        data[301]=154;
        data[300]=153;
        data[299]=152;
        data[298]=152;
        data[297]=151;
        data[296]=151;
        data[295]=150;
        data[294]=150;
        data[293]=149;
        data[292]=149;
        data[291]=148;
        data[290]=148;
        data[289]=147;
        data[288]=147;
        data[287]=146;
        data[286]=146;
        data[285]=145;
        data[284]=145;
        data[283]=144;
        data[282]=144;
        data[281]=143;
        data[280]=143;
        data[279]=142;
        data[278]=142;
        data[277]=141;
        data[276]=141;
        data[275]=140;
        data[274]=140;
        data[273]=139;
        data[272]=139;
        data[271]=138;
        data[270]=138;
        data[269]=137;
        data[268]=137;
        data[267]=136;
        data[266]=136;
        data[265]=135;
        data[264]=135;
        data[263]=134;
        data[262]=134;
        data[261]=133;
        data[260]=133;
        data[259]=132;
        data[258]=132;
        data[257]=131;
        data[256]=131;
        data[255]=130;
        data[254]=130;
        data[253]=129;
        data[252]=129;
        data[251]=128;
        data[250]=128;
        data[249]=127;
        data[248]=126;
        data[247]=126;
        data[246]=125;
        data[245]=125;
        data[244]=124;
        data[243]=124;
        data[242]=123;
        data[241]=123;
        data[240]=122;
        data[239]=122;
        data[238]=121;
        data[237]=121;
        data[236]=120;
        data[235]=120;
        data[234]=119;
        data[233]=119;
        data[232]=118;
        data[231]=118;
        data[230]=117;
        data[229]=117;
        data[228]=116;
        data[227]=116;
        data[226]=115;
        data[225]=115;
        data[224]=114;
        data[223]=114;
        data[222]=113;
        data[221]=113;
        data[220]=112;
        data[219]=112;
        data[218]=111;
        data[217]=111;
        data[216]=110;
        data[215]=110;
        data[214]=109;
        data[213]=109;
        data[212]=108;
        data[211]=108;
        data[210]=107;
        data[209]=107;
        data[208]=106;
        data[207]=106;
        data[206]=105;
        data[205]=105;
        data[204]=104;
        data[203]=104;
        data[202]=103;
        data[201]=103;
        data[200]=102;
        data[199]=101;
        data[198]=101;
        data[197]=100;
        data[196]=100;
        data[195]=99;
        data[194]=99;
        data[193]=98;
        data[192]=98;
        data[191]=97;
        data[190]=97;
        data[189]=96;
        data[188]=96;
        data[187]=95;
        data[186]=95;
        data[185]=94;
        data[184]=94;
        data[183]=93;
        data[182]=93;
        data[181]=92;
        data[180]=92;
        data[179]=91;
        data[178]=91;
        data[177]=90;
        data[176]=90;
        data[175]=89;
        data[174]=89;
        data[173]=88;
        data[172]=88;
        data[171]=87;
        data[170]=87;
        data[169]=86;
        data[168]=86;
        data[167]=85;
        data[166]=85;
        data[165]=84;
        data[164]=84;
        data[163]=83;
        data[162]=83;
        data[161]=82;
        data[160]=82;
        data[159]=81;
        data[158]=81;
        data[157]=80;
        data[156]=80;
        data[155]=79;
        data[154]=79;
        data[153]=78;
        data[152]=78;
        data[151]=77;
        data[150]=77;
        data[149]=76;
        data[148]=75;
        data[147]=75;
        data[146]=74;
        data[145]=74;
        data[144]=73;
        data[143]=73;
        data[142]=72;
        data[141]=72;
        data[140]=71;
        data[139]=71;
        data[138]=70;
        data[137]=70;
        data[136]=69;
        data[135]=69;
        data[134]=68;
        data[133]=68;
        data[132]=67;
        data[131]=67;
        data[130]=66;
        data[129]=66;
        data[128]=65;
        data[127]=65;
        data[126]=64;
        data[125]=64;
        data[124]=63;
        data[123]=63;
        data[122]=62;
        data[121]=62;
        data[120]=61;
        data[119]=61;
        data[118]=60;
        data[117]=60;
        data[116]=59;
        data[115]=59;
        data[114]=58;
        data[113]=58;
        data[112]=57;
        data[111]=57;
        data[110]=56;
        data[109]=56;
        data[108]=55;
        data[107]=55;
        data[106]=54;
        data[105]=54;
        data[104]=53;
        data[103]=53;
        data[102]=52;
        data[101]=52;
        data[100]=51;
        data[99]=50;
        data[98]=50;
        data[97]=49;
        data[96]=49;
        data[95]=48;
        data[94]=48;
        data[93]=47;
        data[92]=47;
        data[91]=46;
        data[90]=46;
        data[89]=45;
        data[88]=45;
        data[87]=44;
        data[86]=44;
        data[85]=43;
        data[84]=43;
        data[83]=42;
        data[82]=42;
        data[81]=41;
        data[80]=41;
        data[79]=40;
        data[78]=40;
        data[77]=39;
        data[76]=39;
        data[75]=38;
        data[74]=38;
        data[73]=37;
        data[72]=37;
        data[71]=36;
        data[70]=36;
        data[69]=35;
        data[68]=35;
        data[67]=34;
        data[66]=34;
        data[65]=33;
        data[64]=33;
        data[63]=32;
        data[62]=32;
        data[61]=31;
        data[60]=31;
        data[59]=30;
        data[58]=30;
        data[57]=29;
        data[56]=29;
        data[55]=28;
        data[54]=28;
        data[53]=27;
        data[52]=27;
        data[51]=26;
        data[50]=25;
        data[49]=25;
        data[48]=24;
        data[47]=24;
        data[46]=23;
        data[45]=23;
        data[44]=22;
        data[43]=22;
        data[42]=21;
        data[41]=21;
        data[40]=20;
        data[39]=20;
        data[38]=19;
        data[37]=19;
        data[36]=18;
        data[35]=18;
        data[34]=17;
        data[33]=17;
        data[32]=16;
        data[31]=16;
        data[30]=15;
        data[29]=15;
        data[28]=14;
        data[27]=14;
        data[26]=13;
        data[25]=13;
        data[24]=12;
        data[23]=12;
        data[22]=11;
        data[21]=11;
        data[20]=10;
        data[19]=10;
        data[18]=9;
        data[17]=9;
        data[16]=8;
        data[15]=8;
        data[14]=7;
        data[13]=7;
        data[12]=6;
        data[11]=6;
        data[10]=5;
        data[9]=5;
        data[8]=4;
        data[7]=4;
        data[6]=3;
        data[5]=3;
        data[4]=2;
        data[3]=2;
        data[2]=1;
        data[1]=1;
        data[0]=0;

    end
     always @(posedge clk) begin
        otp<=data[count];
        count<=(count+1'b1)%mod;
    end
endmodule