module romtatal (
    clk,
    choose,
    cout,
    otp
);
    input clk;
    input [1:0] choose;
    output reg[7:0] otp;
    output reg cout;
    reg [7:0] data[4095:0];
    reg [9:0] count;
    reg [9:0] mod;
   
    initial begin
        cout=0;
         otp=0;
         count=0;
        mod=1000;
        data[4095]=255;
        data[4094]=255;
        data[4093]=255;
        data[4092]=255;
        data[4091]=255;
        data[4090]=255;
        data[4089]=255;
        data[4088]=255;
        data[4087]=255;
        data[4086]=255;
        data[4085]=255;
        data[4084]=255;
        data[4083]=255;
        data[4082]=255;
        data[4081]=255;
        data[4080]=255;
        data[4079]=255;
        data[4078]=255;
        data[4077]=255;
        data[4076]=255;
        data[4075]=255;
        data[4074]=255;
        data[4073]=255;
        data[4072]=255;
        data[4071]=255;
        data[4070]=252;
        data[4069]=250;
        data[4068]=247;
        data[4067]=245;
        data[4066]=242;
        data[4065]=240;
        data[4064]=237;
        data[4063]=235;
        data[4062]=232;
        data[4061]=230;
        data[4060]=227;
        data[4059]=224;
        data[4058]=222;
        data[4057]=219;
        data[4056]=217;
        data[4055]=214;
        data[4054]=212;
        data[4053]=209;
        data[4052]=207;
        data[4051]=204;
        data[4050]=201;
        data[4049]=199;
        data[4048]=196;
        data[4047]=194;
        data[4046]=191;
        data[4045]=189;
        data[4044]=186;
        data[4043]=184;
        data[4042]=181;
        data[4041]=178;
        data[4040]=176;
        data[4039]=173;
        data[4038]=171;
        data[4037]=168;
        data[4036]=166;
        data[4035]=163;
        data[4034]=161;
        data[4033]=158;
        data[4032]=156;
        data[4031]=153;
        data[4030]=150;
        data[4029]=148;
        data[4028]=145;
        data[4027]=143;
        data[4026]=140;
        data[4025]=138;
        data[4024]=135;
        data[4023]=133;
        data[4022]=130;
        data[4021]=128;
        data[4020]=125;
        data[4019]=122;
        data[4018]=120;
        data[4017]=117;
        data[4016]=115;
        data[4015]=112;
        data[4014]=110;
        data[4013]=107;
        data[4012]=105;
        data[4011]=102;
        data[4010]=99;
        data[4009]=97;
        data[4008]=94;
        data[4007]=92;
        data[4006]=89;
        data[4005]=87;
        data[4004]=84;
        data[4003]=82;
        data[4002]=79;
        data[4001]=76;
        data[4000]=74;
        data[3999]=71;
        data[3998]=69;
        data[3997]=66;
        data[3996]=64;
        data[3995]=61;
        data[3994]=59;
        data[3993]=56;
        data[3992]=54;
        data[3991]=51;
        data[3990]=48;
        data[3989]=46;
        data[3988]=43;
        data[3987]=41;
        data[3986]=38;
        data[3985]=36;
        data[3984]=33;
        data[3983]=31;
        data[3982]=28;
        data[3981]=26;
        data[3980]=23;
        data[3979]=20;
        data[3978]=18;
        data[3977]=15;
        data[3976]=13;
        data[3975]=10;
        data[3974]=8;
        data[3973]=5;
        data[3972]=3;
        data[3971]=0;
        data[3970]=1;
        data[3969]=1;
        data[3968]=1;
        data[3967]=1;
        data[3966]=2;
        data[3965]=2;
        data[3964]=2;
        data[3963]=3;
        data[3962]=3;
        data[3961]=3;
        data[3960]=3;
        data[3959]=4;
        data[3958]=4;
        data[3957]=4;
        data[3956]=5;
        data[3955]=5;
        data[3954]=5;
        data[3953]=5;
        data[3952]=6;
        data[3951]=6;
        data[3950]=6;
        data[3949]=7;
        data[3948]=7;
        data[3947]=7;
        data[3946]=7;
        data[3945]=8;
        data[3944]=8;
        data[3943]=8;
        data[3942]=8;
        data[3941]=9;
        data[3940]=9;
        data[3939]=9;
        data[3938]=10;
        data[3937]=10;
        data[3936]=10;
        data[3935]=10;
        data[3934]=11;
        data[3933]=11;
        data[3932]=11;
        data[3931]=12;
        data[3930]=12;
        data[3929]=12;
        data[3928]=12;
        data[3927]=13;
        data[3926]=13;
        data[3925]=13;
        data[3924]=14;
        data[3923]=14;
        data[3922]=14;
        data[3921]=14;
        data[3920]=15;
        data[3919]=15;
        data[3918]=15;
        data[3917]=16;
        data[3916]=16;
        data[3915]=16;
        data[3914]=16;
        data[3913]=17;
        data[3912]=17;
        data[3911]=17;
        data[3910]=18;
        data[3909]=18;
        data[3908]=18;
        data[3907]=18;
        data[3906]=19;
        data[3905]=19;
        data[3904]=19;
        data[3903]=20;
        data[3902]=20;
        data[3901]=20;
        data[3900]=20;
        data[3899]=21;
        data[3898]=21;
        data[3897]=21;
        data[3896]=22;
        data[3895]=22;
        data[3894]=22;
        data[3893]=22;
        data[3892]=23;
        data[3891]=23;
        data[3890]=23;
        data[3889]=24;
        data[3888]=24;
        data[3887]=24;
        data[3886]=24;
        data[3885]=25;
        data[3884]=25;
        data[3883]=25;
        data[3882]=26;
        data[3881]=26;
        data[3880]=26;
        data[3879]=26;
        data[3878]=27;
        data[3877]=27;
        data[3876]=27;
        data[3875]=27;
        data[3874]=28;
        data[3873]=28;
        data[3872]=28;
        data[3871]=29;
        data[3870]=29;
        data[3869]=29;
        data[3868]=29;
        data[3867]=30;
        data[3866]=30;
        data[3865]=30;
        data[3864]=31;
        data[3863]=31;
        data[3862]=31;
        data[3861]=31;
        data[3860]=32;
        data[3859]=32;
        data[3858]=32;
        data[3857]=33;
        data[3856]=33;
        data[3855]=33;
        data[3854]=33;
        data[3853]=34;
        data[3852]=34;
        data[3851]=34;
        data[3850]=35;
        data[3849]=35;
        data[3848]=35;
        data[3847]=35;
        data[3846]=36;
        data[3845]=36;
        data[3844]=36;
        data[3843]=37;
        data[3842]=37;
        data[3841]=37;
        data[3840]=37;
        data[3839]=38;
        data[3838]=38;
        data[3837]=38;
        data[3836]=39;
        data[3835]=39;
        data[3834]=39;
        data[3833]=39;
        data[3832]=40;
        data[3831]=40;
        data[3830]=40;
        data[3829]=41;
        data[3828]=41;
        data[3827]=41;
        data[3826]=41;
        data[3825]=42;
        data[3824]=42;
        data[3823]=42;
        data[3822]=42;
        data[3821]=43;
        data[3820]=43;
        data[3819]=43;
        data[3818]=44;
        data[3817]=44;
        data[3816]=44;
        data[3815]=44;
        data[3814]=45;
        data[3813]=45;
        data[3812]=45;
        data[3811]=46;
        data[3810]=46;
        data[3809]=46;
        data[3808]=46;
        data[3807]=47;
        data[3806]=47;
        data[3805]=47;
        data[3804]=48;
        data[3803]=48;
        data[3802]=48;
        data[3801]=48;
        data[3800]=49;
        data[3799]=49;
        data[3798]=49;
        data[3797]=50;
        data[3796]=50;
        data[3795]=50;
        data[3794]=50;
        data[3793]=51;
        data[3792]=51;
        data[3791]=51;
        data[3790]=52;
        data[3789]=52;
        data[3788]=52;
        data[3787]=52;
        data[3786]=53;
        data[3785]=53;
        data[3784]=53;
        data[3783]=54;
        data[3782]=54;
        data[3781]=54;
        data[3780]=54;
        data[3779]=55;
        data[3778]=55;
        data[3777]=55;
        data[3776]=56;
        data[3775]=56;
        data[3774]=56;
        data[3773]=56;
        data[3772]=57;
        data[3771]=57;
        data[3770]=57;
        data[3769]=58;
        data[3768]=58;
        data[3767]=58;
        data[3766]=58;
        data[3765]=59;
        data[3764]=59;
        data[3763]=59;
        data[3762]=60;
        data[3761]=60;
        data[3760]=60;
        data[3759]=60;
        data[3758]=61;
        data[3757]=61;
        data[3756]=61;
        data[3755]=61;
        data[3754]=62;
        data[3753]=62;
        data[3752]=62;
        data[3751]=63;
        data[3750]=63;
        data[3749]=63;
        data[3748]=63;
        data[3747]=64;
        data[3746]=64;
        data[3745]=64;
        data[3744]=65;
        data[3743]=65;
        data[3742]=65;
        data[3741]=65;
        data[3740]=66;
        data[3739]=66;
        data[3738]=66;
        data[3737]=67;
        data[3736]=67;
        data[3735]=67;
        data[3734]=67;
        data[3733]=68;
        data[3732]=68;
        data[3731]=68;
        data[3730]=69;
        data[3729]=69;
        data[3728]=69;
        data[3727]=69;
        data[3726]=70;
        data[3725]=70;
        data[3724]=70;
        data[3723]=71;
        data[3722]=71;
        data[3721]=71;
        data[3720]=71;
        data[3719]=72;
        data[3718]=72;
        data[3717]=72;
        data[3716]=73;
        data[3715]=73;
        data[3714]=73;
        data[3713]=73;
        data[3712]=74;
        data[3711]=74;
        data[3710]=74;
        data[3709]=75;
        data[3708]=75;
        data[3707]=75;
        data[3706]=75;
        data[3705]=76;
        data[3704]=76;
        data[3703]=76;
        data[3702]=77;
        data[3701]=77;
        data[3700]=77;
        data[3699]=77;
        data[3698]=78;
        data[3697]=78;
        data[3696]=78;
        data[3695]=78;
        data[3694]=79;
        data[3693]=79;
        data[3692]=79;
        data[3691]=80;
        data[3690]=80;
        data[3689]=80;
        data[3688]=80;
        data[3687]=81;
        data[3686]=81;
        data[3685]=81;
        data[3684]=82;
        data[3683]=82;
        data[3682]=82;
        data[3681]=82;
        data[3680]=83;
        data[3679]=83;
        data[3678]=83;
        data[3677]=84;
        data[3676]=84;
        data[3675]=84;
        data[3674]=84;
        data[3673]=85;
        data[3672]=85;
        data[3671]=85;
        data[3670]=86;
        data[3669]=86;
        data[3668]=86;
        data[3667]=86;
        data[3666]=87;
        data[3665]=87;
        data[3664]=87;
        data[3663]=88;
        data[3662]=88;
        data[3661]=88;
        data[3660]=88;
        data[3659]=89;
        data[3658]=89;
        data[3657]=89;
        data[3656]=90;
        data[3655]=90;
        data[3654]=90;
        data[3653]=90;
        data[3652]=91;
        data[3651]=91;
        data[3650]=91;
        data[3649]=92;
        data[3648]=92;
        data[3647]=92;
        data[3646]=92;
        data[3645]=93;
        data[3644]=93;
        data[3643]=93;
        data[3642]=93;
        data[3641]=94;
        data[3640]=94;
        data[3639]=94;
        data[3638]=95;
        data[3637]=95;
        data[3636]=95;
        data[3635]=95;
        data[3634]=96;
        data[3633]=96;
        data[3632]=96;
        data[3631]=97;
        data[3630]=97;
        data[3629]=97;
        data[3628]=97;
        data[3627]=98;
        data[3626]=98;
        data[3625]=98;
        data[3624]=99;
        data[3623]=99;
        data[3622]=99;
        data[3621]=99;
        data[3620]=100;
        data[3619]=100;
        data[3618]=100;
        data[3617]=101;
        data[3616]=101;
        data[3615]=101;
        data[3614]=101;
        data[3613]=102;
        data[3612]=102;
        data[3611]=102;
        data[3610]=103;
        data[3609]=103;
        data[3608]=103;
        data[3607]=103;
        data[3606]=104;
        data[3605]=104;
        data[3604]=104;
        data[3603]=105;
        data[3602]=105;
        data[3601]=105;
        data[3600]=105;
        data[3599]=106;
        data[3598]=106;
        data[3597]=106;
        data[3596]=107;
        data[3595]=107;
        data[3594]=107;
        data[3593]=107;
        data[3592]=108;
        data[3591]=108;
        data[3590]=108;
        data[3589]=109;
        data[3588]=109;
        data[3587]=109;
        data[3586]=109;
        data[3585]=110;
        data[3584]=110;
        data[3583]=110;
        data[3582]=111;
        data[3581]=111;
        data[3580]=111;
        data[3579]=111;
        data[3578]=112;
        data[3577]=112;
        data[3576]=112;
        data[3575]=112;
        data[3574]=113;
        data[3573]=113;
        data[3572]=113;
        data[3571]=114;
        data[3570]=114;
        data[3569]=114;
        data[3568]=114;
        data[3567]=115;
        data[3566]=115;
        data[3565]=115;
        data[3564]=116;
        data[3563]=116;
        data[3562]=116;
        data[3561]=116;
        data[3560]=117;
        data[3559]=117;
        data[3558]=117;
        data[3557]=118;
        data[3556]=118;
        data[3555]=118;
        data[3554]=118;
        data[3553]=119;
        data[3552]=119;
        data[3551]=119;
        data[3550]=120;
        data[3549]=120;
        data[3548]=120;
        data[3547]=120;
        data[3546]=121;
        data[3545]=121;
        data[3544]=121;
        data[3543]=122;
        data[3542]=122;
        data[3541]=122;
        data[3540]=122;
        data[3539]=123;
        data[3538]=123;
        data[3537]=123;
        data[3536]=124;
        data[3535]=124;
        data[3534]=124;
        data[3533]=124;
        data[3532]=125;
        data[3531]=125;
        data[3530]=125;
        data[3529]=126;
        data[3528]=126;
        data[3527]=126;
        data[3526]=126;
        data[3525]=127;
        data[3524]=127;
        data[3523]=127;
        data[3522]=127;
        data[3521]=128;
        data[3520]=128;
        data[3519]=128;
        data[3518]=129;
        data[3517]=129;
        data[3516]=129;
        data[3515]=129;
        data[3514]=130;
        data[3513]=130;
        data[3512]=130;
        data[3511]=131;
        data[3510]=131;
        data[3509]=131;
        data[3508]=131;
        data[3507]=132;
        data[3506]=132;
        data[3505]=132;
        data[3504]=133;
        data[3503]=133;
        data[3502]=133;
        data[3501]=133;
        data[3500]=134;
        data[3499]=134;
        data[3498]=134;
        data[3497]=135;
        data[3496]=135;
        data[3495]=135;
        data[3494]=135;
        data[3493]=136;
        data[3492]=136;
        data[3491]=136;
        data[3490]=137;
        data[3489]=137;
        data[3488]=137;
        data[3487]=137;
        data[3486]=138;
        data[3485]=138;
        data[3484]=138;
        data[3483]=139;
        data[3482]=139;
        data[3481]=139;
        data[3480]=139;
        data[3479]=140;
        data[3478]=140;
        data[3477]=140;
        data[3476]=141;
        data[3475]=141;
        data[3474]=141;
        data[3473]=141;
        data[3472]=142;
        data[3471]=142;
        data[3470]=142;
        data[3469]=143;
        data[3468]=143;
        data[3467]=143;
        data[3466]=143;
        data[3465]=144;
        data[3464]=144;
        data[3463]=144;
        data[3462]=145;
        data[3461]=145;
        data[3460]=145;
        data[3459]=145;
        data[3458]=146;
        data[3457]=146;
        data[3456]=146;
        data[3455]=146;
        data[3454]=147;
        data[3453]=147;
        data[3452]=147;
        data[3451]=148;
        data[3450]=148;
        data[3449]=148;
        data[3448]=148;
        data[3447]=149;
        data[3446]=149;
        data[3445]=149;
        data[3444]=150;
        data[3443]=150;
        data[3442]=150;
        data[3441]=150;
        data[3440]=151;
        data[3439]=151;
        data[3438]=151;
        data[3437]=152;
        data[3436]=152;
        data[3435]=152;
        data[3434]=152;
        data[3433]=153;
        data[3432]=153;
        data[3431]=153;
        data[3430]=154;
        data[3429]=154;
        data[3428]=154;
        data[3427]=154;
        data[3426]=155;
        data[3425]=155;
        data[3424]=155;
        data[3423]=156;
        data[3422]=156;
        data[3421]=156;
        data[3420]=156;
        data[3419]=157;
        data[3418]=157;
        data[3417]=157;
        data[3416]=158;
        data[3415]=158;
        data[3414]=158;
        data[3413]=158;
        data[3412]=159;
        data[3411]=159;
        data[3410]=159;
        data[3409]=160;
        data[3408]=160;
        data[3407]=160;
        data[3406]=160;
        data[3405]=161;
        data[3404]=161;
        data[3403]=161;
        data[3402]=161;
        data[3401]=162;
        data[3400]=162;
        data[3399]=162;
        data[3398]=163;
        data[3397]=163;
        data[3396]=163;
        data[3395]=163;
        data[3394]=164;
        data[3393]=164;
        data[3392]=164;
        data[3391]=165;
        data[3390]=165;
        data[3389]=165;
        data[3388]=165;
        data[3387]=166;
        data[3386]=166;
        data[3385]=166;
        data[3384]=167;
        data[3383]=167;
        data[3382]=167;
        data[3381]=167;
        data[3380]=168;
        data[3379]=168;
        data[3378]=168;
        data[3377]=169;
        data[3376]=169;
        data[3375]=169;
        data[3374]=169;
        data[3373]=170;
        data[3372]=170;
        data[3371]=170;
        data[3370]=171;
        data[3369]=171;
        data[3368]=171;
        data[3367]=171;
        data[3366]=172;
        data[3365]=172;
        data[3364]=172;
        data[3363]=173;
        data[3362]=173;
        data[3361]=173;
        data[3360]=173;
        data[3359]=174;
        data[3358]=174;
        data[3357]=174;
        data[3356]=175;
        data[3355]=175;
        data[3354]=175;
        data[3353]=175;
        data[3352]=176;
        data[3351]=176;
        data[3350]=176;
        data[3349]=177;
        data[3348]=177;
        data[3347]=177;
        data[3346]=177;
        data[3345]=178;
        data[3344]=178;
        data[3343]=178;
        data[3342]=178;
        data[3341]=179;
        data[3340]=179;
        data[3339]=179;
        data[3338]=180;
        data[3337]=180;
        data[3336]=180;
        data[3335]=180;
        data[3334]=181;
        data[3333]=181;
        data[3332]=181;
        data[3331]=182;
        data[3330]=182;
        data[3329]=182;
        data[3328]=182;
        data[3327]=183;
        data[3326]=183;
        data[3325]=183;
        data[3324]=184;
        data[3323]=184;
        data[3322]=184;
        data[3321]=184;
        data[3320]=185;
        data[3319]=185;
        data[3318]=185;
        data[3317]=186;
        data[3316]=186;
        data[3315]=186;
        data[3314]=186;
        data[3313]=187;
        data[3312]=187;
        data[3311]=187;
        data[3310]=188;
        data[3309]=188;
        data[3308]=188;
        data[3307]=188;
        data[3306]=189;
        data[3305]=189;
        data[3304]=189;
        data[3303]=190;
        data[3302]=190;
        data[3301]=190;
        data[3300]=190;
        data[3299]=191;
        data[3298]=191;
        data[3297]=191;
        data[3296]=192;
        data[3295]=192;
        data[3294]=192;
        data[3293]=192;
        data[3292]=193;
        data[3291]=193;
        data[3290]=193;
        data[3289]=194;
        data[3288]=194;
        data[3287]=194;
        data[3286]=194;
        data[3285]=195;
        data[3284]=195;
        data[3283]=195;
        data[3282]=196;
        data[3281]=196;
        data[3280]=196;
        data[3279]=196;
        data[3278]=197;
        data[3277]=197;
        data[3276]=197;
        data[3275]=197;
        data[3274]=198;
        data[3273]=198;
        data[3272]=198;
        data[3271]=199;
        data[3270]=199;
        data[3269]=199;
        data[3268]=199;
        data[3267]=200;
        data[3266]=200;
        data[3265]=200;
        data[3264]=201;
        data[3263]=201;
        data[3262]=201;
        data[3261]=201;
        data[3260]=202;
        data[3259]=202;
        data[3258]=202;
        data[3257]=203;
        data[3256]=203;
        data[3255]=203;
        data[3254]=203;
        data[3253]=204;
        data[3252]=204;
        data[3251]=204;
        data[3250]=205;
        data[3249]=205;
        data[3248]=205;
        data[3247]=205;
        data[3246]=206;
        data[3245]=206;
        data[3244]=206;
        data[3243]=207;
        data[3242]=207;
        data[3241]=207;
        data[3240]=207;
        data[3239]=208;
        data[3238]=208;
        data[3237]=208;
        data[3236]=209;
        data[3235]=209;
        data[3234]=209;
        data[3233]=209;
        data[3232]=210;
        data[3231]=210;
        data[3230]=210;
        data[3229]=211;
        data[3228]=211;
        data[3227]=211;
        data[3226]=211;
        data[3225]=212;
        data[3224]=212;
        data[3223]=212;
        data[3222]=212;
        data[3221]=213;
        data[3220]=213;
        data[3219]=213;
        data[3218]=214;
        data[3217]=214;
        data[3216]=214;
        data[3215]=214;
        data[3214]=215;
        data[3213]=215;
        data[3212]=215;
        data[3211]=216;
        data[3210]=216;
        data[3209]=216;
        data[3208]=216;
        data[3207]=217;
        data[3206]=217;
        data[3205]=217;
        data[3204]=218;
        data[3203]=218;
        data[3202]=218;
        data[3201]=218;
        data[3200]=219;
        data[3199]=219;
        data[3198]=219;
        data[3197]=220;
        data[3196]=220;
        data[3195]=220;
        data[3194]=220;
        data[3193]=221;
        data[3192]=221;
        data[3191]=221;
        data[3190]=222;
        data[3189]=222;
        data[3188]=222;
        data[3187]=222;
        data[3186]=223;
        data[3185]=223;
        data[3184]=223;
        data[3183]=224;
        data[3182]=224;
        data[3181]=224;
        data[3180]=224;
        data[3179]=225;
        data[3178]=225;
        data[3177]=225;
        data[3176]=226;
        data[3175]=226;
        data[3174]=226;
        data[3173]=226;
        data[3172]=227;
        data[3171]=227;
        data[3170]=227;
        data[3169]=228;
        data[3168]=228;
        data[3167]=228;
        data[3166]=228;
        data[3165]=229;
        data[3164]=229;
        data[3163]=229;
        data[3162]=230;
        data[3161]=230;
        data[3160]=230;
        data[3159]=230;
        data[3158]=231;
        data[3157]=231;
        data[3156]=231;
        data[3155]=231;
        data[3154]=232;
        data[3153]=232;
        data[3152]=232;
        data[3151]=233;
        data[3150]=233;
        data[3149]=233;
        data[3148]=233;
        data[3147]=234;
        data[3146]=234;
        data[3145]=234;
        data[3144]=235;
        data[3143]=235;
        data[3142]=235;
        data[3141]=235;
        data[3140]=236;
        data[3139]=236;
        data[3138]=236;
        data[3137]=237;
        data[3136]=237;
        data[3135]=237;
        data[3134]=237;
        data[3133]=238;
        data[3132]=238;
        data[3131]=238;
        data[3130]=239;
        data[3129]=239;
        data[3128]=239;
        data[3127]=239;
        data[3126]=240;
        data[3125]=240;
        data[3124]=240;
        data[3123]=241;
        data[3122]=241;
        data[3121]=241;
        data[3120]=241;
        data[3119]=242;
        data[3118]=242;
        data[3117]=242;
        data[3116]=243;
        data[3115]=243;
        data[3114]=243;
        data[3113]=243;
        data[3112]=244;
        data[3111]=244;
        data[3110]=244;
        data[3109]=245;
        data[3108]=245;
        data[3107]=245;
        data[3106]=245;
        data[3105]=246;
        data[3104]=246;
        data[3103]=246;
        data[3102]=246;
        data[3101]=247;
        data[3100]=247;
        data[3099]=247;
        data[3098]=248;
        data[3097]=248;
        data[3096]=248;
        data[3095]=248;
        data[3094]=249;
        data[3093]=249;
        data[3092]=249;
        data[3091]=250;
        data[3090]=250;
        data[3089]=250;
        data[3088]=250;
        data[3087]=251;
        data[3086]=251;
        data[3085]=251;
        data[3084]=252;
        data[3083]=252;
        data[3082]=252;
        data[3081]=252;
        data[3080]=253;
        data[3079]=253;
        data[3078]=253;
        data[3077]=254;
        data[3076]=254;
        data[3075]=254;
        data[3074]=254;
        data[3073]=255;
        data[3072]=255;
        data[3071]=255;
        data[3070]=255;
        data[3069]=255;
        data[3068]=255;
        data[3067]=255;
        data[3066]=255;
        data[3065]=255;
        data[3064]=255;
        data[3063]=255;
        data[3062]=255;
        data[3061]=255;
        data[3060]=255;
        data[3059]=255;
        data[3058]=255;
        data[3057]=255;
        data[3056]=255;
        data[3055]=255;
        data[3054]=255;
        data[3053]=255;
        data[3052]=255;
        data[3051]=255;
        data[3050]=255;
        data[3049]=255;
        data[3048]=255;
        data[3047]=255;
        data[3046]=254;
        data[3045]=254;
        data[3044]=253;
        data[3043]=253;
        data[3042]=252;
        data[3041]=252;
        data[3040]=251;
        data[3039]=251;
        data[3038]=250;
        data[3037]=250;
        data[3036]=249;
        data[3035]=249;
        data[3034]=248;
        data[3033]=248;
        data[3032]=247;
        data[3031]=247;
        data[3030]=246;
        data[3029]=246;
        data[3028]=245;
        data[3027]=245;
        data[3026]=244;
        data[3025]=244;
        data[3024]=243;
        data[3023]=243;
        data[3022]=242;
        data[3021]=242;
        data[3020]=241;
        data[3019]=241;
        data[3018]=240;
        data[3017]=240;
        data[3016]=239;
        data[3015]=239;
        data[3014]=238;
        data[3013]=238;
        data[3012]=237;
        data[3011]=237;
        data[3010]=236;
        data[3009]=236;
        data[3008]=235;
        data[3007]=235;
        data[3006]=234;
        data[3005]=234;
        data[3004]=233;
        data[3003]=233;
        data[3002]=232;
        data[3001]=232;
        data[3000]=231;
        data[2999]=231;
        data[2998]=230;
        data[2997]=230;
        data[2996]=229;
        data[2995]=228;
        data[2994]=228;
        data[2993]=227;
        data[2992]=227;
        data[2991]=226;
        data[2990]=226;
        data[2989]=225;
        data[2988]=225;
        data[2987]=224;
        data[2986]=224;
        data[2985]=223;
        data[2984]=223;
        data[2983]=222;
        data[2982]=222;
        data[2981]=221;
        data[2980]=221;
        data[2979]=220;
        data[2978]=220;
        data[2977]=219;
        data[2976]=219;
        data[2975]=218;
        data[2974]=218;
        data[2973]=217;
        data[2972]=217;
        data[2971]=216;
        data[2970]=216;
        data[2969]=215;
        data[2968]=215;
        data[2967]=214;
        data[2966]=214;
        data[2965]=213;
        data[2964]=213;
        data[2963]=212;
        data[2962]=212;
        data[2961]=211;
        data[2960]=211;
        data[2959]=210;
        data[2958]=210;
        data[2957]=209;
        data[2956]=209;
        data[2955]=208;
        data[2954]=208;
        data[2953]=207;
        data[2952]=207;
        data[2951]=206;
        data[2950]=206;
        data[2949]=205;
        data[2948]=205;
        data[2947]=204;
        data[2946]=203;
        data[2945]=203;
        data[2944]=202;
        data[2943]=202;
        data[2942]=201;
        data[2941]=201;
        data[2940]=200;
        data[2939]=200;
        data[2938]=199;
        data[2937]=199;
        data[2936]=198;
        data[2935]=198;
        data[2934]=197;
        data[2933]=197;
        data[2932]=196;
        data[2931]=196;
        data[2930]=195;
        data[2929]=195;
        data[2928]=194;
        data[2927]=194;
        data[2926]=193;
        data[2925]=193;
        data[2924]=192;
        data[2923]=192;
        data[2922]=191;
        data[2921]=191;
        data[2920]=190;
        data[2919]=190;
        data[2918]=189;
        data[2917]=189;
        data[2916]=188;
        data[2915]=188;
        data[2914]=187;
        data[2913]=187;
        data[2912]=186;
        data[2911]=186;
        data[2910]=185;
        data[2909]=185;
        data[2908]=184;
        data[2907]=184;
        data[2906]=183;
        data[2905]=183;
        data[2904]=182;
        data[2903]=182;
        data[2902]=181;
        data[2901]=181;
        data[2900]=180;
        data[2899]=180;
        data[2898]=179;
        data[2897]=178;
        data[2896]=178;
        data[2895]=177;
        data[2894]=177;
        data[2893]=176;
        data[2892]=176;
        data[2891]=175;
        data[2890]=175;
        data[2889]=174;
        data[2888]=174;
        data[2887]=173;
        data[2886]=173;
        data[2885]=172;
        data[2884]=172;
        data[2883]=171;
        data[2882]=171;
        data[2881]=170;
        data[2880]=170;
        data[2879]=169;
        data[2878]=169;
        data[2877]=168;
        data[2876]=168;
        data[2875]=167;
        data[2874]=167;
        data[2873]=166;
        data[2872]=166;
        data[2871]=165;
        data[2870]=165;
        data[2869]=164;
        data[2868]=164;
        data[2867]=163;
        data[2866]=163;
        data[2865]=162;
        data[2864]=162;
        data[2863]=161;
        data[2862]=161;
        data[2861]=160;
        data[2860]=160;
        data[2859]=159;
        data[2858]=159;
        data[2857]=158;
        data[2856]=158;
        data[2855]=157;
        data[2854]=157;
        data[2853]=156;
        data[2852]=156;
        data[2851]=155;
        data[2850]=155;
        data[2849]=154;
        data[2848]=154;
        data[2847]=153;
        data[2846]=152;
        data[2845]=152;
        data[2844]=151;
        data[2843]=151;
        data[2842]=150;
        data[2841]=150;
        data[2840]=149;
        data[2839]=149;
        data[2838]=148;
        data[2837]=148;
        data[2836]=147;
        data[2835]=147;
        data[2834]=146;
        data[2833]=146;
        data[2832]=145;
        data[2831]=145;
        data[2830]=144;
        data[2829]=144;
        data[2828]=143;
        data[2827]=143;
        data[2826]=142;
        data[2825]=142;
        data[2824]=141;
        data[2823]=141;
        data[2822]=140;
        data[2821]=140;
        data[2820]=139;
        data[2819]=139;
        data[2818]=138;
        data[2817]=138;
        data[2816]=137;
        data[2815]=137;
        data[2814]=136;
        data[2813]=136;
        data[2812]=135;
        data[2811]=135;
        data[2810]=134;
        data[2809]=134;
        data[2808]=133;
        data[2807]=133;
        data[2806]=132;
        data[2805]=132;
        data[2804]=131;
        data[2803]=131;
        data[2802]=130;
        data[2801]=130;
        data[2800]=129;
        data[2799]=129;
        data[2798]=128;
        data[2797]=127;
        data[2796]=127;
        data[2795]=126;
        data[2794]=126;
        data[2793]=125;
        data[2792]=125;
        data[2791]=124;
        data[2790]=124;
        data[2789]=123;
        data[2788]=123;
        data[2787]=122;
        data[2786]=122;
        data[2785]=121;
        data[2784]=121;
        data[2783]=120;
        data[2782]=120;
        data[2781]=119;
        data[2780]=119;
        data[2779]=118;
        data[2778]=118;
        data[2777]=117;
        data[2776]=117;
        data[2775]=116;
        data[2774]=116;
        data[2773]=115;
        data[2772]=115;
        data[2771]=114;
        data[2770]=114;
        data[2769]=113;
        data[2768]=113;
        data[2767]=112;
        data[2766]=112;
        data[2765]=111;
        data[2764]=111;
        data[2763]=110;
        data[2762]=110;
        data[2761]=109;
        data[2760]=109;
        data[2759]=108;
        data[2758]=108;
        data[2757]=107;
        data[2756]=107;
        data[2755]=106;
        data[2754]=106;
        data[2753]=105;
        data[2752]=105;
        data[2751]=104;
        data[2750]=104;
        data[2749]=103;
        data[2748]=103;
        data[2747]=102;
        data[2746]=101;
        data[2745]=101;
        data[2744]=100;
        data[2743]=100;
        data[2742]=99;
        data[2741]=99;
        data[2740]=98;
        data[2739]=98;
        data[2738]=97;
        data[2737]=97;
        data[2736]=96;
        data[2735]=96;
        data[2734]=95;
        data[2733]=95;
        data[2732]=94;
        data[2731]=94;
        data[2730]=93;
        data[2729]=93;
        data[2728]=92;
        data[2727]=92;
        data[2726]=91;
        data[2725]=91;
        data[2724]=90;
        data[2723]=90;
        data[2722]=89;
        data[2721]=89;
        data[2720]=88;
        data[2719]=88;
        data[2718]=87;
        data[2717]=87;
        data[2716]=86;
        data[2715]=86;
        data[2714]=85;
        data[2713]=85;
        data[2712]=84;
        data[2711]=84;
        data[2710]=83;
        data[2709]=83;
        data[2708]=82;
        data[2707]=82;
        data[2706]=81;
        data[2705]=81;
        data[2704]=80;
        data[2703]=80;
        data[2702]=79;
        data[2701]=79;
        data[2700]=78;
        data[2699]=78;
        data[2698]=77;
        data[2697]=76;
        data[2696]=76;
        data[2695]=75;
        data[2694]=75;
        data[2693]=74;
        data[2692]=74;
        data[2691]=73;
        data[2690]=73;
        data[2689]=72;
        data[2688]=72;
        data[2687]=71;
        data[2686]=71;
        data[2685]=70;
        data[2684]=70;
        data[2683]=69;
        data[2682]=69;
        data[2681]=68;
        data[2680]=68;
        data[2679]=67;
        data[2678]=67;
        data[2677]=66;
        data[2676]=66;
        data[2675]=65;
        data[2674]=65;
        data[2673]=64;
        data[2672]=64;
        data[2671]=63;
        data[2670]=63;
        data[2669]=62;
        data[2668]=62;
        data[2667]=61;
        data[2666]=61;
        data[2665]=60;
        data[2664]=60;
        data[2663]=59;
        data[2662]=59;
        data[2661]=58;
        data[2660]=58;
        data[2659]=57;
        data[2658]=57;
        data[2657]=56;
        data[2656]=56;
        data[2655]=55;
        data[2654]=55;
        data[2653]=54;
        data[2652]=54;
        data[2651]=53;
        data[2650]=53;
        data[2649]=52;
        data[2648]=52;
        data[2647]=51;
        data[2646]=50;
        data[2645]=50;
        data[2644]=49;
        data[2643]=49;
        data[2642]=48;
        data[2641]=48;
        data[2640]=47;
        data[2639]=47;
        data[2638]=46;
        data[2637]=46;
        data[2636]=45;
        data[2635]=45;
        data[2634]=44;
        data[2633]=44;
        data[2632]=43;
        data[2631]=43;
        data[2630]=42;
        data[2629]=42;
        data[2628]=41;
        data[2627]=41;
        data[2626]=40;
        data[2625]=40;
        data[2624]=39;
        data[2623]=39;
        data[2622]=38;
        data[2621]=38;
        data[2620]=37;
        data[2619]=37;
        data[2618]=36;
        data[2617]=36;
        data[2616]=35;
        data[2615]=35;
        data[2614]=34;
        data[2613]=34;
        data[2612]=33;
        data[2611]=33;
        data[2610]=32;
        data[2609]=32;
        data[2608]=31;
        data[2607]=31;
        data[2606]=30;
        data[2605]=30;
        data[2604]=29;
        data[2603]=29;
        data[2602]=28;
        data[2601]=28;
        data[2600]=27;
        data[2599]=27;
        data[2598]=26;
        data[2597]=25;
        data[2596]=25;
        data[2595]=24;
        data[2594]=24;
        data[2593]=23;
        data[2592]=23;
        data[2591]=22;
        data[2590]=22;
        data[2589]=21;
        data[2588]=21;
        data[2587]=20;
        data[2586]=20;
        data[2585]=19;
        data[2584]=19;
        data[2583]=18;
        data[2582]=18;
        data[2581]=17;
        data[2580]=17;
        data[2579]=16;
        data[2578]=16;
        data[2577]=15;
        data[2576]=15;
        data[2575]=14;
        data[2574]=14;
        data[2573]=13;
        data[2572]=13;
        data[2571]=12;
        data[2570]=12;
        data[2569]=11;
        data[2568]=11;
        data[2567]=10;
        data[2566]=10;
        data[2565]=9;
        data[2564]=9;
        data[2563]=8;
        data[2562]=8;
        data[2561]=7;
        data[2560]=7;
        data[2559]=6;
        data[2558]=6;
        data[2557]=5;
        data[2556]=5;
        data[2555]=4;
        data[2554]=4;
        data[2553]=3;
        data[2552]=3;
        data[2551]=2;
        data[2550]=2;
        data[2549]=1;
        data[2548]=1;
        data[2547]=1;
        data[2546]=1;
        data[2545]=2;
        data[2544]=2;
        data[2543]=3;
        data[2542]=3;
        data[2541]=4;
        data[2540]=4;
        data[2539]=5;
        data[2538]=5;
        data[2537]=6;
        data[2536]=6;
        data[2535]=7;
        data[2534]=7;
        data[2533]=8;
        data[2532]=8;
        data[2531]=9;
        data[2530]=9;
        data[2529]=10;
        data[2528]=10;
        data[2527]=11;
        data[2526]=11;
        data[2525]=12;
        data[2524]=12;
        data[2523]=13;
        data[2522]=13;
        data[2521]=14;
        data[2520]=14;
        data[2519]=15;
        data[2518]=15;
        data[2517]=16;
        data[2516]=16;
        data[2515]=17;
        data[2514]=17;
        data[2513]=18;
        data[2512]=18;
        data[2511]=19;
        data[2510]=19;
        data[2509]=20;
        data[2508]=20;
        data[2507]=21;
        data[2506]=21;
        data[2505]=22;
        data[2504]=22;
        data[2503]=23;
        data[2502]=23;
        data[2501]=24;
        data[2500]=24;
        data[2499]=25;
        data[2498]=25;
        data[2497]=26;
        data[2496]=27;
        data[2495]=27;
        data[2494]=28;
        data[2493]=28;
        data[2492]=29;
        data[2491]=29;
        data[2490]=30;
        data[2489]=30;
        data[2488]=31;
        data[2487]=31;
        data[2486]=32;
        data[2485]=32;
        data[2484]=33;
        data[2483]=33;
        data[2482]=34;
        data[2481]=34;
        data[2480]=35;
        data[2479]=35;
        data[2478]=36;
        data[2477]=36;
        data[2476]=37;
        data[2475]=37;
        data[2474]=38;
        data[2473]=38;
        data[2472]=39;
        data[2471]=39;
        data[2470]=40;
        data[2469]=40;
        data[2468]=41;
        data[2467]=41;
        data[2466]=42;
        data[2465]=42;
        data[2464]=43;
        data[2463]=43;
        data[2462]=44;
        data[2461]=44;
        data[2460]=45;
        data[2459]=45;
        data[2458]=46;
        data[2457]=46;
        data[2456]=47;
        data[2455]=47;
        data[2454]=48;
        data[2453]=48;
        data[2452]=49;
        data[2451]=49;
        data[2450]=50;
        data[2449]=50;
        data[2448]=51;
        data[2447]=52;
        data[2446]=52;
        data[2445]=53;
        data[2444]=53;
        data[2443]=54;
        data[2442]=54;
        data[2441]=55;
        data[2440]=55;
        data[2439]=56;
        data[2438]=56;
        data[2437]=57;
        data[2436]=57;
        data[2435]=58;
        data[2434]=58;
        data[2433]=59;
        data[2432]=59;
        data[2431]=60;
        data[2430]=60;
        data[2429]=61;
        data[2428]=61;
        data[2427]=62;
        data[2426]=62;
        data[2425]=63;
        data[2424]=63;
        data[2423]=64;
        data[2422]=64;
        data[2421]=65;
        data[2420]=65;
        data[2419]=66;
        data[2418]=66;
        data[2417]=67;
        data[2416]=67;
        data[2415]=68;
        data[2414]=68;
        data[2413]=69;
        data[2412]=69;
        data[2411]=70;
        data[2410]=70;
        data[2409]=71;
        data[2408]=71;
        data[2407]=72;
        data[2406]=72;
        data[2405]=73;
        data[2404]=73;
        data[2403]=74;
        data[2402]=74;
        data[2401]=75;
        data[2400]=75;
        data[2399]=76;
        data[2398]=76;
        data[2397]=77;
        data[2396]=78;
        data[2395]=78;
        data[2394]=79;
        data[2393]=79;
        data[2392]=80;
        data[2391]=80;
        data[2390]=81;
        data[2389]=81;
        data[2388]=82;
        data[2387]=82;
        data[2386]=83;
        data[2385]=83;
        data[2384]=84;
        data[2383]=84;
        data[2382]=85;
        data[2381]=85;
        data[2380]=86;
        data[2379]=86;
        data[2378]=87;
        data[2377]=87;
        data[2376]=88;
        data[2375]=88;
        data[2374]=89;
        data[2373]=89;
        data[2372]=90;
        data[2371]=90;
        data[2370]=91;
        data[2369]=91;
        data[2368]=92;
        data[2367]=92;
        data[2366]=93;
        data[2365]=93;
        data[2364]=94;
        data[2363]=94;
        data[2362]=95;
        data[2361]=95;
        data[2360]=96;
        data[2359]=96;
        data[2358]=97;
        data[2357]=97;
        data[2356]=98;
        data[2355]=98;
        data[2354]=99;
        data[2353]=99;
        data[2352]=100;
        data[2351]=100;
        data[2350]=101;
        data[2349]=101;
        data[2348]=102;
        data[2347]=103;
        data[2346]=103;
        data[2345]=104;
        data[2344]=104;
        data[2343]=105;
        data[2342]=105;
        data[2341]=106;
        data[2340]=106;
        data[2339]=107;
        data[2338]=107;
        data[2337]=108;
        data[2336]=108;
        data[2335]=109;
        data[2334]=109;
        data[2333]=110;
        data[2332]=110;
        data[2331]=111;
        data[2330]=111;
        data[2329]=112;
        data[2328]=112;
        data[2327]=113;
        data[2326]=113;
        data[2325]=114;
        data[2324]=114;
        data[2323]=115;
        data[2322]=115;
        data[2321]=116;
        data[2320]=116;
        data[2319]=117;
        data[2318]=117;
        data[2317]=118;
        data[2316]=118;
        data[2315]=119;
        data[2314]=119;
        data[2313]=120;
        data[2312]=120;
        data[2311]=121;
        data[2310]=121;
        data[2309]=122;
        data[2308]=122;
        data[2307]=123;
        data[2306]=123;
        data[2305]=124;
        data[2304]=124;
        data[2303]=125;
        data[2302]=125;
        data[2301]=126;
        data[2300]=126;
        data[2299]=127;
        data[2298]=127;
        data[2297]=128;
        data[2296]=129;
        data[2295]=129;
        data[2294]=130;
        data[2293]=130;
        data[2292]=131;
        data[2291]=131;
        data[2290]=132;
        data[2289]=132;
        data[2288]=133;
        data[2287]=133;
        data[2286]=134;
        data[2285]=134;
        data[2284]=135;
        data[2283]=135;
        data[2282]=136;
        data[2281]=136;
        data[2280]=137;
        data[2279]=137;
        data[2278]=138;
        data[2277]=138;
        data[2276]=139;
        data[2275]=139;
        data[2274]=140;
        data[2273]=140;
        data[2272]=141;
        data[2271]=141;
        data[2270]=142;
        data[2269]=142;
        data[2268]=143;
        data[2267]=143;
        data[2266]=144;
        data[2265]=144;
        data[2264]=145;
        data[2263]=145;
        data[2262]=146;
        data[2261]=146;
        data[2260]=147;
        data[2259]=147;
        data[2258]=148;
        data[2257]=148;
        data[2256]=149;
        data[2255]=149;
        data[2254]=150;
        data[2253]=150;
        data[2252]=151;
        data[2251]=151;
        data[2250]=152;
        data[2249]=152;
        data[2248]=153;
        data[2247]=154;
        data[2246]=154;
        data[2245]=155;
        data[2244]=155;
        data[2243]=156;
        data[2242]=156;
        data[2241]=157;
        data[2240]=157;
        data[2239]=158;
        data[2238]=158;
        data[2237]=159;
        data[2236]=159;
        data[2235]=160;
        data[2234]=160;
        data[2233]=161;
        data[2232]=161;
        data[2231]=162;
        data[2230]=162;
        data[2229]=163;
        data[2228]=163;
        data[2227]=164;
        data[2226]=164;
        data[2225]=165;
        data[2224]=165;
        data[2223]=166;
        data[2222]=166;
        data[2221]=167;
        data[2220]=167;
        data[2219]=168;
        data[2218]=168;
        data[2217]=169;
        data[2216]=169;
        data[2215]=170;
        data[2214]=170;
        data[2213]=171;
        data[2212]=171;
        data[2211]=172;
        data[2210]=172;
        data[2209]=173;
        data[2208]=173;
        data[2207]=174;
        data[2206]=174;
        data[2205]=175;
        data[2204]=175;
        data[2203]=176;
        data[2202]=176;
        data[2201]=177;
        data[2200]=177;
        data[2199]=178;
        data[2198]=178;
        data[2197]=179;
        data[2196]=180;
        data[2195]=180;
        data[2194]=181;
        data[2193]=181;
        data[2192]=182;
        data[2191]=182;
        data[2190]=183;
        data[2189]=183;
        data[2188]=184;
        data[2187]=184;
        data[2186]=185;
        data[2185]=185;
        data[2184]=186;
        data[2183]=186;
        data[2182]=187;
        data[2181]=187;
        data[2180]=188;
        data[2179]=188;
        data[2178]=189;
        data[2177]=189;
        data[2176]=190;
        data[2175]=190;
        data[2174]=191;
        data[2173]=191;
        data[2172]=192;
        data[2171]=192;
        data[2170]=193;
        data[2169]=193;
        data[2168]=194;
        data[2167]=194;
        data[2166]=195;
        data[2165]=195;
        data[2164]=196;
        data[2163]=196;
        data[2162]=197;
        data[2161]=197;
        data[2160]=198;
        data[2159]=198;
        data[2158]=199;
        data[2157]=199;
        data[2156]=200;
        data[2155]=200;
        data[2154]=201;
        data[2153]=201;
        data[2152]=202;
        data[2151]=202;
        data[2150]=203;
        data[2149]=203;
        data[2148]=204;
        data[2147]=205;
        data[2146]=205;
        data[2145]=206;
        data[2144]=206;
        data[2143]=207;
        data[2142]=207;
        data[2141]=208;
        data[2140]=208;
        data[2139]=209;
        data[2138]=209;
        data[2137]=210;
        data[2136]=210;
        data[2135]=211;
        data[2134]=211;
        data[2133]=212;
        data[2132]=212;
        data[2131]=213;
        data[2130]=213;
        data[2129]=214;
        data[2128]=214;
        data[2127]=215;
        data[2126]=215;
        data[2125]=216;
        data[2124]=216;
        data[2123]=217;
        data[2122]=217;
        data[2121]=218;
        data[2120]=218;
        data[2119]=219;
        data[2118]=219;
        data[2117]=220;
        data[2116]=220;
        data[2115]=221;
        data[2114]=221;
        data[2113]=222;
        data[2112]=222;
        data[2111]=223;
        data[2110]=223;
        data[2109]=224;
        data[2108]=224;
        data[2107]=225;
        data[2106]=225;
        data[2105]=226;
        data[2104]=226;
        data[2103]=227;
        data[2102]=227;
        data[2101]=228;
        data[2100]=228;
        data[2099]=229;
        data[2098]=230;
        data[2097]=230;
        data[2096]=231;
        data[2095]=231;
        data[2094]=232;
        data[2093]=232;
        data[2092]=233;
        data[2091]=233;
        data[2090]=234;
        data[2089]=234;
        data[2088]=235;
        data[2087]=235;
        data[2086]=236;
        data[2085]=236;
        data[2084]=237;
        data[2083]=237;
        data[2082]=238;
        data[2081]=238;
        data[2080]=239;
        data[2079]=239;
        data[2078]=240;
        data[2077]=240;
        data[2076]=241;
        data[2075]=241;
        data[2074]=242;
        data[2073]=242;
        data[2072]=243;
        data[2071]=243;
        data[2070]=244;
        data[2069]=244;
        data[2068]=245;
        data[2067]=245;
        data[2066]=246;
        data[2065]=246;
        data[2064]=247;
        data[2063]=247;
        data[2062]=248;
        data[2061]=248;
        data[2060]=249;
        data[2059]=249;
        data[2058]=250;
        data[2057]=250;
        data[2056]=251;
        data[2055]=251;
        data[2054]=252;
        data[2053]=252;
        data[2052]=253;
        data[2051]=253;
        data[2050]=254;
        data[2049]=254;
        data[2048]=255;
        data[2047]=255;
        data[2046]=255;
        data[2045]=255;
        data[2044]=255;
        data[2043]=255;
        data[2042]=255;
        data[2041]=255;
        data[2040]=255;
        data[2039]=255;
        data[2038]=255;
        data[2037]=255;
        data[2036]=255;
        data[2035]=255;
        data[2034]=255;
        data[2033]=255;
        data[2032]=255;
        data[2031]=255;
        data[2030]=255;
        data[2029]=255;
        data[2028]=255;
        data[2027]=255;
        data[2026]=255;
        data[2025]=255;
        data[2024]=255;
        data[2023]=0;
        data[2022]=0;
        data[2021]=0;
        data[2020]=0;
        data[2019]=0;
        data[2018]=0;
        data[2017]=0;
        data[2016]=0;
        data[2015]=0;
        data[2014]=0;
        data[2013]=0;
        data[2012]=0;
        data[2011]=0;
        data[2010]=0;
        data[2009]=0;
        data[2008]=0;
        data[2007]=0;
        data[2006]=0;
        data[2005]=0;
        data[2004]=0;
        data[2003]=0;
        data[2002]=0;
        data[2001]=0;
        data[2000]=0;
        data[1999]=0;
        data[1998]=0;
        data[1997]=0;
        data[1996]=0;
        data[1995]=0;
        data[1994]=0;
        data[1993]=0;
        data[1992]=0;
        data[1991]=0;
        data[1990]=0;
        data[1989]=0;
        data[1988]=0;
        data[1987]=0;
        data[1986]=0;
        data[1985]=0;
        data[1984]=0;
        data[1983]=0;
        data[1982]=0;
        data[1981]=0;
        data[1980]=0;
        data[1979]=0;
        data[1978]=0;
        data[1977]=0;
        data[1976]=0;
        data[1975]=0;
        data[1974]=0;
        data[1973]=0;
        data[1972]=0;
        data[1971]=0;
        data[1970]=0;
        data[1969]=0;
        data[1968]=0;
        data[1967]=0;
        data[1966]=0;
        data[1965]=0;
        data[1964]=0;
        data[1963]=0;
        data[1962]=0;
        data[1961]=0;
        data[1960]=0;
        data[1959]=0;
        data[1958]=0;
        data[1957]=0;
        data[1956]=0;
        data[1955]=0;
        data[1954]=0;
        data[1953]=0;
        data[1952]=0;
        data[1951]=0;
        data[1950]=0;
        data[1949]=0;
        data[1948]=0;
        data[1947]=0;
        data[1946]=0;
        data[1945]=0;
        data[1944]=0;
        data[1943]=0;
        data[1942]=0;
        data[1941]=0;
        data[1940]=0;
        data[1939]=0;
        data[1938]=0;
        data[1937]=0;
        data[1936]=0;
        data[1935]=0;
        data[1934]=0;
        data[1933]=0;
        data[1932]=0;
        data[1931]=0;
        data[1930]=0;
        data[1929]=0;
        data[1928]=0;
        data[1927]=0;
        data[1926]=0;
        data[1925]=0;
        data[1924]=0;
        data[1923]=0;
        data[1922]=0;
        data[1921]=0;
        data[1920]=0;
        data[1919]=0;
        data[1918]=0;
        data[1917]=0;
        data[1916]=0;
        data[1915]=0;
        data[1914]=0;
        data[1913]=0;
        data[1912]=0;
        data[1911]=0;
        data[1910]=0;
        data[1909]=0;
        data[1908]=0;
        data[1907]=0;
        data[1906]=0;
        data[1905]=0;
        data[1904]=0;
        data[1903]=0;
        data[1902]=0;
        data[1901]=0;
        data[1900]=0;
        data[1899]=0;
        data[1898]=0;
        data[1897]=0;
        data[1896]=0;
        data[1895]=0;
        data[1894]=0;
        data[1893]=0;
        data[1892]=0;
        data[1891]=0;
        data[1890]=0;
        data[1889]=0;
        data[1888]=0;
        data[1887]=0;
        data[1886]=0;
        data[1885]=0;
        data[1884]=0;
        data[1883]=0;
        data[1882]=0;
        data[1881]=0;
        data[1880]=0;
        data[1879]=0;
        data[1878]=0;
        data[1877]=0;
        data[1876]=0;
        data[1875]=0;
        data[1874]=0;
        data[1873]=0;
        data[1872]=0;
        data[1871]=0;
        data[1870]=0;
        data[1869]=0;
        data[1868]=0;
        data[1867]=0;
        data[1866]=0;
        data[1865]=0;
        data[1864]=0;
        data[1863]=0;
        data[1862]=0;
        data[1861]=0;
        data[1860]=0;
        data[1859]=0;
        data[1858]=0;
        data[1857]=0;
        data[1856]=0;
        data[1855]=0;
        data[1854]=0;
        data[1853]=0;
        data[1852]=0;
        data[1851]=0;
        data[1850]=0;
        data[1849]=0;
        data[1848]=0;
        data[1847]=0;
        data[1846]=0;
        data[1845]=0;
        data[1844]=0;
        data[1843]=0;
        data[1842]=0;
        data[1841]=0;
        data[1840]=0;
        data[1839]=0;
        data[1838]=0;
        data[1837]=0;
        data[1836]=0;
        data[1835]=0;
        data[1834]=0;
        data[1833]=0;
        data[1832]=0;
        data[1831]=0;
        data[1830]=0;
        data[1829]=0;
        data[1828]=0;
        data[1827]=0;
        data[1826]=0;
        data[1825]=0;
        data[1824]=0;
        data[1823]=0;
        data[1822]=0;
        data[1821]=0;
        data[1820]=0;
        data[1819]=0;
        data[1818]=0;
        data[1817]=0;
        data[1816]=0;
        data[1815]=0;
        data[1814]=0;
        data[1813]=0;
        data[1812]=0;
        data[1811]=0;
        data[1810]=0;
        data[1809]=0;
        data[1808]=0;
        data[1807]=0;
        data[1806]=0;
        data[1805]=0;
        data[1804]=0;
        data[1803]=0;
        data[1802]=0;
        data[1801]=0;
        data[1800]=0;
        data[1799]=0;
        data[1798]=0;
        data[1797]=0;
        data[1796]=0;
        data[1795]=0;
        data[1794]=0;
        data[1793]=0;
        data[1792]=0;
        data[1791]=0;
        data[1790]=0;
        data[1789]=0;
        data[1788]=0;
        data[1787]=0;
        data[1786]=0;
        data[1785]=0;
        data[1784]=0;
        data[1783]=0;
        data[1782]=0;
        data[1781]=0;
        data[1780]=0;
        data[1779]=0;
        data[1778]=0;
        data[1777]=0;
        data[1776]=0;
        data[1775]=0;
        data[1774]=0;
        data[1773]=0;
        data[1772]=0;
        data[1771]=0;
        data[1770]=0;
        data[1769]=0;
        data[1768]=0;
        data[1767]=0;
        data[1766]=0;
        data[1765]=0;
        data[1764]=0;
        data[1763]=0;
        data[1762]=0;
        data[1761]=0;
        data[1760]=0;
        data[1759]=0;
        data[1758]=0;
        data[1757]=0;
        data[1756]=0;
        data[1755]=0;
        data[1754]=0;
        data[1753]=0;
        data[1752]=0;
        data[1751]=0;
        data[1750]=0;
        data[1749]=0;
        data[1748]=0;
        data[1747]=0;
        data[1746]=0;
        data[1745]=0;
        data[1744]=0;
        data[1743]=0;
        data[1742]=0;
        data[1741]=0;
        data[1740]=0;
        data[1739]=0;
        data[1738]=0;
        data[1737]=0;
        data[1736]=0;
        data[1735]=0;
        data[1734]=0;
        data[1733]=0;
        data[1732]=0;
        data[1731]=0;
        data[1730]=0;
        data[1729]=0;
        data[1728]=0;
        data[1727]=0;
        data[1726]=0;
        data[1725]=0;
        data[1724]=0;
        data[1723]=0;
        data[1722]=0;
        data[1721]=0;
        data[1720]=0;
        data[1719]=0;
        data[1718]=0;
        data[1717]=0;
        data[1716]=0;
        data[1715]=0;
        data[1714]=0;
        data[1713]=0;
        data[1712]=0;
        data[1711]=0;
        data[1710]=0;
        data[1709]=0;
        data[1708]=0;
        data[1707]=0;
        data[1706]=0;
        data[1705]=0;
        data[1704]=0;
        data[1703]=0;
        data[1702]=0;
        data[1701]=0;
        data[1700]=0;
        data[1699]=0;
        data[1698]=0;
        data[1697]=0;
        data[1696]=0;
        data[1695]=0;
        data[1694]=0;
        data[1693]=0;
        data[1692]=0;
        data[1691]=0;
        data[1690]=0;
        data[1689]=0;
        data[1688]=0;
        data[1687]=0;
        data[1686]=0;
        data[1685]=0;
        data[1684]=0;
        data[1683]=0;
        data[1682]=0;
        data[1681]=0;
        data[1680]=0;
        data[1679]=0;
        data[1678]=0;
        data[1677]=0;
        data[1676]=0;
        data[1675]=0;
        data[1674]=0;
        data[1673]=0;
        data[1672]=0;
        data[1671]=0;
        data[1670]=0;
        data[1669]=0;
        data[1668]=0;
        data[1667]=0;
        data[1666]=0;
        data[1665]=0;
        data[1664]=0;
        data[1663]=0;
        data[1662]=0;
        data[1661]=0;
        data[1660]=0;
        data[1659]=0;
        data[1658]=0;
        data[1657]=0;
        data[1656]=0;
        data[1655]=0;
        data[1654]=0;
        data[1653]=0;
        data[1652]=0;
        data[1651]=0;
        data[1650]=0;
        data[1649]=0;
        data[1648]=0;
        data[1647]=0;
        data[1646]=0;
        data[1645]=0;
        data[1644]=0;
        data[1643]=0;
        data[1642]=0;
        data[1641]=0;
        data[1640]=0;
        data[1639]=0;
        data[1638]=0;
        data[1637]=0;
        data[1636]=0;
        data[1635]=0;
        data[1634]=0;
        data[1633]=0;
        data[1632]=0;
        data[1631]=0;
        data[1630]=0;
        data[1629]=0;
        data[1628]=0;
        data[1627]=0;
        data[1626]=0;
        data[1625]=0;
        data[1624]=0;
        data[1623]=0;
        data[1622]=0;
        data[1621]=0;
        data[1620]=0;
        data[1619]=0;
        data[1618]=0;
        data[1617]=0;
        data[1616]=0;
        data[1615]=0;
        data[1614]=0;
        data[1613]=0;
        data[1612]=0;
        data[1611]=0;
        data[1610]=0;
        data[1609]=0;
        data[1608]=0;
        data[1607]=0;
        data[1606]=0;
        data[1605]=0;
        data[1604]=0;
        data[1603]=0;
        data[1602]=0;
        data[1601]=0;
        data[1600]=0;
        data[1599]=0;
        data[1598]=0;
        data[1597]=0;
        data[1596]=0;
        data[1595]=0;
        data[1594]=0;
        data[1593]=0;
        data[1592]=0;
        data[1591]=0;
        data[1590]=0;
        data[1589]=0;
        data[1588]=0;
        data[1587]=0;
        data[1586]=0;
        data[1585]=0;
        data[1584]=0;
        data[1583]=0;
        data[1582]=0;
        data[1581]=0;
        data[1580]=0;
        data[1579]=0;
        data[1578]=0;
        data[1577]=0;
        data[1576]=0;
        data[1575]=0;
        data[1574]=0;
        data[1573]=0;
        data[1572]=0;
        data[1571]=0;
        data[1570]=0;
        data[1569]=0;
        data[1568]=0;
        data[1567]=0;
        data[1566]=0;
        data[1565]=0;
        data[1564]=0;
        data[1563]=0;
        data[1562]=0;
        data[1561]=0;
        data[1560]=0;
        data[1559]=0;
        data[1558]=0;
        data[1557]=0;
        data[1556]=0;
        data[1555]=0;
        data[1554]=0;
        data[1553]=0;
        data[1552]=0;
        data[1551]=0;
        data[1550]=0;
        data[1549]=0;
        data[1548]=0;
        data[1547]=0;
        data[1546]=0;
        data[1545]=0;
        data[1544]=0;
        data[1543]=0;
        data[1542]=0;
        data[1541]=0;
        data[1540]=0;
        data[1539]=0;
        data[1538]=0;
        data[1537]=0;
        data[1536]=0;
        data[1535]=0;
        data[1534]=0;
        data[1533]=0;
        data[1532]=0;
        data[1531]=0;
        data[1530]=0;
        data[1529]=0;
        data[1528]=0;
        data[1527]=0;
        data[1526]=0;
        data[1525]=0;
        data[1524]=0;
        data[1523]=255;
        data[1522]=255;
        data[1521]=255;
        data[1520]=255;
        data[1519]=255;
        data[1518]=255;
        data[1517]=255;
        data[1516]=255;
        data[1515]=255;
        data[1514]=255;
        data[1513]=255;
        data[1512]=255;
        data[1511]=255;
        data[1510]=255;
        data[1509]=255;
        data[1508]=255;
        data[1507]=255;
        data[1506]=255;
        data[1505]=255;
        data[1504]=255;
        data[1503]=255;
        data[1502]=255;
        data[1501]=255;
        data[1500]=255;
        data[1499]=255;
        data[1498]=255;
        data[1497]=255;
        data[1496]=255;
        data[1495]=255;
        data[1494]=255;
        data[1493]=255;
        data[1492]=255;
        data[1491]=255;
        data[1490]=255;
        data[1489]=255;
        data[1488]=255;
        data[1487]=255;
        data[1486]=255;
        data[1485]=255;
        data[1484]=255;
        data[1483]=255;
        data[1482]=255;
        data[1481]=255;
        data[1480]=255;
        data[1479]=255;
        data[1478]=255;
        data[1477]=255;
        data[1476]=255;
        data[1475]=255;
        data[1474]=255;
        data[1473]=255;
        data[1472]=255;
        data[1471]=255;
        data[1470]=255;
        data[1469]=255;
        data[1468]=255;
        data[1467]=255;
        data[1466]=255;
        data[1465]=255;
        data[1464]=255;
        data[1463]=255;
        data[1462]=255;
        data[1461]=255;
        data[1460]=255;
        data[1459]=255;
        data[1458]=255;
        data[1457]=255;
        data[1456]=255;
        data[1455]=255;
        data[1454]=255;
        data[1453]=255;
        data[1452]=255;
        data[1451]=255;
        data[1450]=255;
        data[1449]=255;
        data[1448]=255;
        data[1447]=255;
        data[1446]=255;
        data[1445]=255;
        data[1444]=255;
        data[1443]=255;
        data[1442]=255;
        data[1441]=255;
        data[1440]=255;
        data[1439]=255;
        data[1438]=255;
        data[1437]=255;
        data[1436]=255;
        data[1435]=255;
        data[1434]=255;
        data[1433]=255;
        data[1432]=255;
        data[1431]=255;
        data[1430]=255;
        data[1429]=255;
        data[1428]=255;
        data[1427]=255;
        data[1426]=255;
        data[1425]=255;
        data[1424]=255;
        data[1423]=255;
        data[1422]=255;
        data[1421]=255;
        data[1420]=255;
        data[1419]=255;
        data[1418]=255;
        data[1417]=255;
        data[1416]=255;
        data[1415]=255;
        data[1414]=255;
        data[1413]=255;
        data[1412]=255;
        data[1411]=255;
        data[1410]=255;
        data[1409]=255;
        data[1408]=255;
        data[1407]=255;
        data[1406]=255;
        data[1405]=255;
        data[1404]=255;
        data[1403]=255;
        data[1402]=255;
        data[1401]=255;
        data[1400]=255;
        data[1399]=255;
        data[1398]=255;
        data[1397]=255;
        data[1396]=255;
        data[1395]=255;
        data[1394]=255;
        data[1393]=255;
        data[1392]=255;
        data[1391]=255;
        data[1390]=255;
        data[1389]=255;
        data[1388]=255;
        data[1387]=255;
        data[1386]=255;
        data[1385]=255;
        data[1384]=255;
        data[1383]=255;
        data[1382]=255;
        data[1381]=255;
        data[1380]=255;
        data[1379]=255;
        data[1378]=255;
        data[1377]=255;
        data[1376]=255;
        data[1375]=255;
        data[1374]=255;
        data[1373]=255;
        data[1372]=255;
        data[1371]=255;
        data[1370]=255;
        data[1369]=255;
        data[1368]=255;
        data[1367]=255;
        data[1366]=255;
        data[1365]=255;
        data[1364]=255;
        data[1363]=255;
        data[1362]=255;
        data[1361]=255;
        data[1360]=255;
        data[1359]=255;
        data[1358]=255;
        data[1357]=255;
        data[1356]=255;
        data[1355]=255;
        data[1354]=255;
        data[1353]=255;
        data[1352]=255;
        data[1351]=255;
        data[1350]=255;
        data[1349]=255;
        data[1348]=255;
        data[1347]=255;
        data[1346]=255;
        data[1345]=255;
        data[1344]=255;
        data[1343]=255;
        data[1342]=255;
        data[1341]=255;
        data[1340]=255;
        data[1339]=255;
        data[1338]=255;
        data[1337]=255;
        data[1336]=255;
        data[1335]=255;
        data[1334]=255;
        data[1333]=255;
        data[1332]=255;
        data[1331]=255;
        data[1330]=255;
        data[1329]=255;
        data[1328]=255;
        data[1327]=255;
        data[1326]=255;
        data[1325]=255;
        data[1324]=255;
        data[1323]=255;
        data[1322]=255;
        data[1321]=255;
        data[1320]=255;
        data[1319]=255;
        data[1318]=255;
        data[1317]=255;
        data[1316]=255;
        data[1315]=255;
        data[1314]=255;
        data[1313]=255;
        data[1312]=255;
        data[1311]=255;
        data[1310]=255;
        data[1309]=255;
        data[1308]=255;
        data[1307]=255;
        data[1306]=255;
        data[1305]=255;
        data[1304]=255;
        data[1303]=255;
        data[1302]=255;
        data[1301]=255;
        data[1300]=255;
        data[1299]=255;
        data[1298]=255;
        data[1297]=255;
        data[1296]=255;
        data[1295]=255;
        data[1294]=255;
        data[1293]=255;
        data[1292]=255;
        data[1291]=255;
        data[1290]=255;
        data[1289]=255;
        data[1288]=255;
        data[1287]=255;
        data[1286]=255;
        data[1285]=255;
        data[1284]=255;
        data[1283]=255;
        data[1282]=255;
        data[1281]=255;
        data[1280]=255;
        data[1279]=255;
        data[1278]=255;
        data[1277]=255;
        data[1276]=255;
        data[1275]=255;
        data[1274]=255;
        data[1273]=255;
        data[1272]=255;
        data[1271]=255;
        data[1270]=255;
        data[1269]=255;
        data[1268]=255;
        data[1267]=255;
        data[1266]=255;
        data[1265]=255;
        data[1264]=255;
        data[1263]=255;
        data[1262]=255;
        data[1261]=255;
        data[1260]=255;
        data[1259]=255;
        data[1258]=255;
        data[1257]=255;
        data[1256]=255;
        data[1255]=255;
        data[1254]=255;
        data[1253]=255;
        data[1252]=255;
        data[1251]=255;
        data[1250]=255;
        data[1249]=255;
        data[1248]=255;
        data[1247]=255;
        data[1246]=255;
        data[1245]=255;
        data[1244]=255;
        data[1243]=255;
        data[1242]=255;
        data[1241]=255;
        data[1240]=255;
        data[1239]=255;
        data[1238]=255;
        data[1237]=255;
        data[1236]=255;
        data[1235]=255;
        data[1234]=255;
        data[1233]=255;
        data[1232]=255;
        data[1231]=255;
        data[1230]=255;
        data[1229]=255;
        data[1228]=255;
        data[1227]=255;
        data[1226]=255;
        data[1225]=255;
        data[1224]=255;
        data[1223]=255;
        data[1222]=255;
        data[1221]=255;
        data[1220]=255;
        data[1219]=255;
        data[1218]=255;
        data[1217]=255;
        data[1216]=255;
        data[1215]=255;
        data[1214]=255;
        data[1213]=255;
        data[1212]=255;
        data[1211]=255;
        data[1210]=255;
        data[1209]=255;
        data[1208]=255;
        data[1207]=255;
        data[1206]=255;
        data[1205]=255;
        data[1204]=255;
        data[1203]=255;
        data[1202]=255;
        data[1201]=255;
        data[1200]=255;
        data[1199]=255;
        data[1198]=255;
        data[1197]=255;
        data[1196]=255;
        data[1195]=255;
        data[1194]=255;
        data[1193]=255;
        data[1192]=255;
        data[1191]=255;
        data[1190]=255;
        data[1189]=255;
        data[1188]=255;
        data[1187]=255;
        data[1186]=255;
        data[1185]=255;
        data[1184]=255;
        data[1183]=255;
        data[1182]=255;
        data[1181]=255;
        data[1180]=255;
        data[1179]=255;
        data[1178]=255;
        data[1177]=255;
        data[1176]=255;
        data[1175]=255;
        data[1174]=255;
        data[1173]=255;
        data[1172]=255;
        data[1171]=255;
        data[1170]=255;
        data[1169]=255;
        data[1168]=255;
        data[1167]=255;
        data[1166]=255;
        data[1165]=255;
        data[1164]=255;
        data[1163]=255;
        data[1162]=255;
        data[1161]=255;
        data[1160]=255;
        data[1159]=255;
        data[1158]=255;
        data[1157]=255;
        data[1156]=255;
        data[1155]=255;
        data[1154]=255;
        data[1153]=255;
        data[1152]=255;
        data[1151]=255;
        data[1150]=255;
        data[1149]=255;
        data[1148]=255;
        data[1147]=255;
        data[1146]=255;
        data[1145]=255;
        data[1144]=255;
        data[1143]=255;
        data[1142]=255;
        data[1141]=255;
        data[1140]=255;
        data[1139]=255;
        data[1138]=255;
        data[1137]=255;
        data[1136]=255;
        data[1135]=255;
        data[1134]=255;
        data[1133]=255;
        data[1132]=255;
        data[1131]=255;
        data[1130]=255;
        data[1129]=255;
        data[1128]=255;
        data[1127]=255;
        data[1126]=255;
        data[1125]=255;
        data[1124]=255;
        data[1123]=255;
        data[1122]=255;
        data[1121]=255;
        data[1120]=255;
        data[1119]=255;
        data[1118]=255;
        data[1117]=255;
        data[1116]=255;
        data[1115]=255;
        data[1114]=255;
        data[1113]=255;
        data[1112]=255;
        data[1111]=255;
        data[1110]=255;
        data[1109]=255;
        data[1108]=255;
        data[1107]=255;
        data[1106]=255;
        data[1105]=255;
        data[1104]=255;
        data[1103]=255;
        data[1102]=255;
        data[1101]=255;
        data[1100]=255;
        data[1099]=255;
        data[1098]=255;
        data[1097]=255;
        data[1096]=255;
        data[1095]=255;
        data[1094]=255;
        data[1093]=255;
        data[1092]=255;
        data[1091]=255;
        data[1090]=255;
        data[1089]=255;
        data[1088]=255;
        data[1087]=255;
        data[1086]=255;
        data[1085]=255;
        data[1084]=255;
        data[1083]=255;
        data[1082]=255;
        data[1081]=255;
        data[1080]=255;
        data[1079]=255;
        data[1078]=255;
        data[1077]=255;
        data[1076]=255;
        data[1075]=255;
        data[1074]=255;
        data[1073]=255;
        data[1072]=255;
        data[1071]=255;
        data[1070]=255;
        data[1069]=255;
        data[1068]=255;
        data[1067]=255;
        data[1066]=255;
        data[1065]=255;
        data[1064]=255;
        data[1063]=255;
        data[1062]=255;
        data[1061]=255;
        data[1060]=255;
        data[1059]=255;
        data[1058]=255;
        data[1057]=255;
        data[1056]=255;
        data[1055]=255;
        data[1054]=255;
        data[1053]=255;
        data[1052]=255;
        data[1051]=255;
        data[1050]=255;
        data[1049]=255;
        data[1048]=255;
        data[1047]=255;
        data[1046]=255;
        data[1045]=255;
        data[1044]=255;
        data[1043]=255;
        data[1042]=255;
        data[1041]=255;
        data[1040]=255;
        data[1039]=255;
        data[1038]=255;
        data[1037]=255;
        data[1036]=255;
        data[1035]=255;
        data[1034]=255;
        data[1033]=255;
        data[1032]=255;
        data[1031]=255;
        data[1030]=255;
        data[1029]=255;
        data[1028]=255;
        data[1027]=255;
        data[1026]=255;
        data[1025]=255;
        data[1024]=255;
        data[1023]=255;
        data[1022]=255;
        data[1021]=255;
        data[1020]=255;
        data[1019]=255;
        data[1018]=255;
        data[1017]=255;
        data[1016]=255;
        data[1015]=255;
        data[1014]=255;
        data[1013]=255;
        data[1012]=255;
        data[1011]=255;
        data[1010]=255;
        data[1009]=255;
        data[1008]=255;
        data[1007]=255;
        data[1006]=255;
        data[1005]=255;
        data[1004]=255;
        data[1003]=255;
        data[1002]=255;
        data[1001]=255;
        data[1000]=255;
        data[999]=129;
        data[998]=130;
        data[997]=130;
        data[996]=131;
        data[995]=132;
        data[994]=133;
        data[993]=134;
        data[992]=134;
        data[991]=135;
        data[990]=136;
        data[989]=137;
        data[988]=138;
        data[987]=138;
        data[986]=139;
        data[985]=140;
        data[984]=141;
        data[983]=142;
        data[982]=142;
        data[981]=143;
        data[980]=144;
        data[979]=145;
        data[978]=146;
        data[977]=146;
        data[976]=147;
        data[975]=148;
        data[974]=149;
        data[973]=150;
        data[972]=150;
        data[971]=151;
        data[970]=152;
        data[969]=153;
        data[968]=154;
        data[967]=154;
        data[966]=155;
        data[965]=156;
        data[964]=157;
        data[963]=157;
        data[962]=158;
        data[961]=159;
        data[960]=160;
        data[959]=161;
        data[958]=161;
        data[957]=162;
        data[956]=163;
        data[955]=164;
        data[954]=164;
        data[953]=165;
        data[952]=166;
        data[951]=167;
        data[950]=168;
        data[949]=168;
        data[948]=169;
        data[947]=170;
        data[946]=171;
        data[945]=171;
        data[944]=172;
        data[943]=173;
        data[942]=174;
        data[941]=174;
        data[940]=175;
        data[939]=176;
        data[938]=177;
        data[937]=177;
        data[936]=178;
        data[935]=179;
        data[934]=180;
        data[933]=180;
        data[932]=181;
        data[931]=182;
        data[930]=182;
        data[929]=183;
        data[928]=184;
        data[927]=185;
        data[926]=185;
        data[925]=186;
        data[924]=187;
        data[923]=188;
        data[922]=188;
        data[921]=189;
        data[920]=190;
        data[919]=190;
        data[918]=191;
        data[917]=192;
        data[916]=192;
        data[915]=193;
        data[914]=194;
        data[913]=195;
        data[912]=195;
        data[911]=196;
        data[910]=197;
        data[909]=197;
        data[908]=198;
        data[907]=199;
        data[906]=199;
        data[905]=200;
        data[904]=201;
        data[903]=201;
        data[902]=202;
        data[901]=203;
        data[900]=203;
        data[899]=204;
        data[898]=205;
        data[897]=205;
        data[896]=206;
        data[895]=206;
        data[894]=207;
        data[893]=208;
        data[892]=208;
        data[891]=209;
        data[890]=210;
        data[889]=210;
        data[888]=211;
        data[887]=211;
        data[886]=212;
        data[885]=213;
        data[884]=213;
        data[883]=214;
        data[882]=214;
        data[881]=215;
        data[880]=216;
        data[879]=216;
        data[878]=217;
        data[877]=217;
        data[876]=218;
        data[875]=219;
        data[874]=219;
        data[873]=220;
        data[872]=220;
        data[871]=221;
        data[870]=221;
        data[869]=222;
        data[868]=222;
        data[867]=223;
        data[866]=223;
        data[865]=224;
        data[864]=225;
        data[863]=225;
        data[862]=226;
        data[861]=226;
        data[860]=227;
        data[859]=227;
        data[858]=228;
        data[857]=228;
        data[856]=229;
        data[855]=229;
        data[854]=230;
        data[853]=230;
        data[852]=231;
        data[851]=231;
        data[850]=232;
        data[849]=232;
        data[848]=232;
        data[847]=233;
        data[846]=233;
        data[845]=234;
        data[844]=234;
        data[843]=235;
        data[842]=235;
        data[841]=236;
        data[840]=236;
        data[839]=237;
        data[838]=237;
        data[837]=237;
        data[836]=238;
        data[835]=238;
        data[834]=239;
        data[833]=239;
        data[832]=239;
        data[831]=240;
        data[830]=240;
        data[829]=241;
        data[828]=241;
        data[827]=241;
        data[826]=242;
        data[825]=242;
        data[824]=242;
        data[823]=243;
        data[822]=243;
        data[821]=243;
        data[820]=244;
        data[819]=244;
        data[818]=244;
        data[817]=245;
        data[816]=245;
        data[815]=245;
        data[814]=246;
        data[813]=246;
        data[812]=246;
        data[811]=247;
        data[810]=247;
        data[809]=247;
        data[808]=248;
        data[807]=248;
        data[806]=248;
        data[805]=248;
        data[804]=249;
        data[803]=249;
        data[802]=249;
        data[801]=249;
        data[800]=250;
        data[799]=250;
        data[798]=250;
        data[797]=250;
        data[796]=251;
        data[795]=251;
        data[794]=251;
        data[793]=251;
        data[792]=252;
        data[791]=252;
        data[790]=252;
        data[789]=252;
        data[788]=252;
        data[787]=253;
        data[786]=253;
        data[785]=253;
        data[784]=253;
        data[783]=253;
        data[782]=253;
        data[781]=254;
        data[780]=254;
        data[779]=254;
        data[778]=254;
        data[777]=254;
        data[776]=254;
        data[775]=254;
        data[774]=255;
        data[773]=255;
        data[772]=255;
        data[771]=255;
        data[770]=255;
        data[769]=255;
        data[768]=255;
        data[767]=255;
        data[766]=255;
        data[765]=255;
        data[764]=255;
        data[763]=255;
        data[762]=255;
        data[761]=255;
        data[760]=255;
        data[759]=255;
        data[758]=255;
        data[757]=255;
        data[756]=255;
        data[755]=255;
        data[754]=255;
        data[753]=255;
        data[752]=255;
        data[751]=255;
        data[750]=255;
        data[749]=255;
        data[748]=255;
        data[747]=255;
        data[746]=255;
        data[745]=255;
        data[744]=255;
        data[743]=255;
        data[742]=255;
        data[741]=255;
        data[740]=255;
        data[739]=255;
        data[738]=255;
        data[737]=255;
        data[736]=255;
        data[735]=255;
        data[734]=255;
        data[733]=255;
        data[732]=255;
        data[731]=255;
        data[730]=255;
        data[729]=255;
        data[728]=255;
        data[727]=255;
        data[726]=255;
        data[725]=254;
        data[724]=254;
        data[723]=254;
        data[722]=254;
        data[721]=254;
        data[720]=254;
        data[719]=254;
        data[718]=253;
        data[717]=253;
        data[716]=253;
        data[715]=253;
        data[714]=253;
        data[713]=253;
        data[712]=252;
        data[711]=252;
        data[710]=252;
        data[709]=252;
        data[708]=252;
        data[707]=251;
        data[706]=251;
        data[705]=251;
        data[704]=251;
        data[703]=250;
        data[702]=250;
        data[701]=250;
        data[700]=250;
        data[699]=249;
        data[698]=249;
        data[697]=249;
        data[696]=249;
        data[695]=248;
        data[694]=248;
        data[693]=248;
        data[692]=248;
        data[691]=247;
        data[690]=247;
        data[689]=247;
        data[688]=246;
        data[687]=246;
        data[686]=246;
        data[685]=245;
        data[684]=245;
        data[683]=245;
        data[682]=244;
        data[681]=244;
        data[680]=244;
        data[679]=243;
        data[678]=243;
        data[677]=243;
        data[676]=242;
        data[675]=242;
        data[674]=242;
        data[673]=241;
        data[672]=241;
        data[671]=241;
        data[670]=240;
        data[669]=240;
        data[668]=239;
        data[667]=239;
        data[666]=239;
        data[665]=238;
        data[664]=238;
        data[663]=237;
        data[662]=237;
        data[661]=237;
        data[660]=236;
        data[659]=236;
        data[658]=235;
        data[657]=235;
        data[656]=234;
        data[655]=234;
        data[654]=233;
        data[653]=233;
        data[652]=232;
        data[651]=232;
        data[650]=232;
        data[649]=231;
        data[648]=231;
        data[647]=230;
        data[646]=230;
        data[645]=229;
        data[644]=229;
        data[643]=228;
        data[642]=228;
        data[641]=227;
        data[640]=227;
        data[639]=226;
        data[638]=226;
        data[637]=225;
        data[636]=225;
        data[635]=224;
        data[634]=223;
        data[633]=223;
        data[632]=222;
        data[631]=222;
        data[630]=221;
        data[629]=221;
        data[628]=220;
        data[627]=220;
        data[626]=219;
        data[625]=219;
        data[624]=218;
        data[623]=217;
        data[622]=217;
        data[621]=216;
        data[620]=216;
        data[619]=215;
        data[618]=214;
        data[617]=214;
        data[616]=213;
        data[615]=213;
        data[614]=212;
        data[613]=211;
        data[612]=211;
        data[611]=210;
        data[610]=210;
        data[609]=209;
        data[608]=208;
        data[607]=208;
        data[606]=207;
        data[605]=206;
        data[604]=206;
        data[603]=205;
        data[602]=205;
        data[601]=204;
        data[600]=203;
        data[599]=203;
        data[598]=202;
        data[597]=201;
        data[596]=201;
        data[595]=200;
        data[594]=199;
        data[593]=199;
        data[592]=198;
        data[591]=197;
        data[590]=197;
        data[589]=196;
        data[588]=195;
        data[587]=195;
        data[586]=194;
        data[585]=193;
        data[584]=192;
        data[583]=192;
        data[582]=191;
        data[581]=190;
        data[580]=190;
        data[579]=189;
        data[578]=188;
        data[577]=188;
        data[576]=187;
        data[575]=186;
        data[574]=185;
        data[573]=185;
        data[572]=184;
        data[571]=183;
        data[570]=182;
        data[569]=182;
        data[568]=181;
        data[567]=180;
        data[566]=180;
        data[565]=179;
        data[564]=178;
        data[563]=177;
        data[562]=177;
        data[561]=176;
        data[560]=175;
        data[559]=174;
        data[558]=174;
        data[557]=173;
        data[556]=172;
        data[555]=171;
        data[554]=171;
        data[553]=170;
        data[552]=169;
        data[551]=168;
        data[550]=168;
        data[549]=167;
        data[548]=166;
        data[547]=165;
        data[546]=164;
        data[545]=164;
        data[544]=163;
        data[543]=162;
        data[542]=161;
        data[541]=161;
        data[540]=160;
        data[539]=159;
        data[538]=158;
        data[537]=157;
        data[536]=157;
        data[535]=156;
        data[534]=155;
        data[533]=154;
        data[532]=154;
        data[531]=153;
        data[530]=152;
        data[529]=151;
        data[528]=150;
        data[527]=150;
        data[526]=149;
        data[525]=148;
        data[524]=147;
        data[523]=146;
        data[522]=146;
        data[521]=145;
        data[520]=144;
        data[519]=143;
        data[518]=142;
        data[517]=142;
        data[516]=141;
        data[515]=140;
        data[514]=139;
        data[513]=138;
        data[512]=138;
        data[511]=137;
        data[510]=136;
        data[509]=135;
        data[508]=134;
        data[507]=134;
        data[506]=133;
        data[505]=132;
        data[504]=131;
        data[503]=130;
        data[502]=130;
        data[501]=129;
        data[500]=128;
        data[499]=127;
        data[498]=126;
        data[497]=126;
        data[496]=125;
        data[495]=124;
        data[494]=123;
        data[493]=122;
        data[492]=122;
        data[491]=121;
        data[490]=120;
        data[489]=119;
        data[488]=118;
        data[487]=118;
        data[486]=117;
        data[485]=116;
        data[484]=115;
        data[483]=114;
        data[482]=114;
        data[481]=113;
        data[480]=112;
        data[479]=111;
        data[478]=110;
        data[477]=110;
        data[476]=109;
        data[475]=108;
        data[474]=107;
        data[473]=106;
        data[472]=106;
        data[471]=105;
        data[470]=104;
        data[469]=103;
        data[468]=102;
        data[467]=102;
        data[466]=101;
        data[465]=100;
        data[464]=99;
        data[463]=99;
        data[462]=98;
        data[461]=97;
        data[460]=96;
        data[459]=95;
        data[458]=95;
        data[457]=94;
        data[456]=93;
        data[455]=92;
        data[454]=92;
        data[453]=91;
        data[452]=90;
        data[451]=89;
        data[450]=88;
        data[449]=88;
        data[448]=87;
        data[447]=86;
        data[446]=85;
        data[445]=85;
        data[444]=84;
        data[443]=83;
        data[442]=82;
        data[441]=82;
        data[440]=81;
        data[439]=80;
        data[438]=79;
        data[437]=79;
        data[436]=78;
        data[435]=77;
        data[434]=76;
        data[433]=76;
        data[432]=75;
        data[431]=74;
        data[430]=74;
        data[429]=73;
        data[428]=72;
        data[427]=71;
        data[426]=71;
        data[425]=70;
        data[424]=69;
        data[423]=68;
        data[422]=68;
        data[421]=67;
        data[420]=66;
        data[419]=66;
        data[418]=65;
        data[417]=64;
        data[416]=64;
        data[415]=63;
        data[414]=62;
        data[413]=61;
        data[412]=61;
        data[411]=60;
        data[410]=59;
        data[409]=59;
        data[408]=58;
        data[407]=57;
        data[406]=57;
        data[405]=56;
        data[404]=55;
        data[403]=55;
        data[402]=54;
        data[401]=53;
        data[400]=53;
        data[399]=52;
        data[398]=51;
        data[397]=51;
        data[396]=50;
        data[395]=50;
        data[394]=49;
        data[393]=48;
        data[392]=48;
        data[391]=47;
        data[390]=46;
        data[389]=46;
        data[388]=45;
        data[387]=45;
        data[386]=44;
        data[385]=43;
        data[384]=43;
        data[383]=42;
        data[382]=42;
        data[381]=41;
        data[380]=40;
        data[379]=40;
        data[378]=39;
        data[377]=39;
        data[376]=38;
        data[375]=37;
        data[374]=37;
        data[373]=36;
        data[372]=36;
        data[371]=35;
        data[370]=35;
        data[369]=34;
        data[368]=34;
        data[367]=33;
        data[366]=33;
        data[365]=32;
        data[364]=31;
        data[363]=31;
        data[362]=30;
        data[361]=30;
        data[360]=29;
        data[359]=29;
        data[358]=28;
        data[357]=28;
        data[356]=27;
        data[355]=27;
        data[354]=26;
        data[353]=26;
        data[352]=25;
        data[351]=25;
        data[350]=24;
        data[349]=24;
        data[348]=24;
        data[347]=23;
        data[346]=23;
        data[345]=22;
        data[344]=22;
        data[343]=21;
        data[342]=21;
        data[341]=20;
        data[340]=20;
        data[339]=19;
        data[338]=19;
        data[337]=19;
        data[336]=18;
        data[335]=18;
        data[334]=17;
        data[333]=17;
        data[332]=17;
        data[331]=16;
        data[330]=16;
        data[329]=15;
        data[328]=15;
        data[327]=15;
        data[326]=14;
        data[325]=14;
        data[324]=14;
        data[323]=13;
        data[322]=13;
        data[321]=13;
        data[320]=12;
        data[319]=12;
        data[318]=12;
        data[317]=11;
        data[316]=11;
        data[315]=11;
        data[314]=10;
        data[313]=10;
        data[312]=10;
        data[311]=9;
        data[310]=9;
        data[309]=9;
        data[308]=8;
        data[307]=8;
        data[306]=8;
        data[305]=8;
        data[304]=7;
        data[303]=7;
        data[302]=7;
        data[301]=7;
        data[300]=6;
        data[299]=6;
        data[298]=6;
        data[297]=6;
        data[296]=5;
        data[295]=5;
        data[294]=5;
        data[293]=5;
        data[292]=4;
        data[291]=4;
        data[290]=4;
        data[289]=4;
        data[288]=4;
        data[287]=3;
        data[286]=3;
        data[285]=3;
        data[284]=3;
        data[283]=3;
        data[282]=3;
        data[281]=2;
        data[280]=2;
        data[279]=2;
        data[278]=2;
        data[277]=2;
        data[276]=2;
        data[275]=2;
        data[274]=1;
        data[273]=1;
        data[272]=1;
        data[271]=1;
        data[270]=1;
        data[269]=1;
        data[268]=1;
        data[267]=1;
        data[266]=1;
        data[265]=1;
        data[264]=0;
        data[263]=0;
        data[262]=0;
        data[261]=0;
        data[260]=0;
        data[259]=0;
        data[258]=0;
        data[257]=0;
        data[256]=0;
        data[255]=0;
        data[254]=0;
        data[253]=0;
        data[252]=0;
        data[251]=0;
        data[250]=0;
        data[249]=0;
        data[248]=0;
        data[247]=0;
        data[246]=0;
        data[245]=0;
        data[244]=0;
        data[243]=0;
        data[242]=0;
        data[241]=0;
        data[240]=0;
        data[239]=0;
        data[238]=0;
        data[237]=0;
        data[236]=0;
        data[235]=1;
        data[234]=1;
        data[233]=1;
        data[232]=1;
        data[231]=1;
        data[230]=1;
        data[229]=1;
        data[228]=1;
        data[227]=1;
        data[226]=1;
        data[225]=2;
        data[224]=2;
        data[223]=2;
        data[222]=2;
        data[221]=2;
        data[220]=2;
        data[219]=2;
        data[218]=3;
        data[217]=3;
        data[216]=3;
        data[215]=3;
        data[214]=3;
        data[213]=3;
        data[212]=4;
        data[211]=4;
        data[210]=4;
        data[209]=4;
        data[208]=4;
        data[207]=5;
        data[206]=5;
        data[205]=5;
        data[204]=5;
        data[203]=6;
        data[202]=6;
        data[201]=6;
        data[200]=6;
        data[199]=7;
        data[198]=7;
        data[197]=7;
        data[196]=7;
        data[195]=8;
        data[194]=8;
        data[193]=8;
        data[192]=8;
        data[191]=9;
        data[190]=9;
        data[189]=9;
        data[188]=10;
        data[187]=10;
        data[186]=10;
        data[185]=11;
        data[184]=11;
        data[183]=11;
        data[182]=12;
        data[181]=12;
        data[180]=12;
        data[179]=13;
        data[178]=13;
        data[177]=13;
        data[176]=14;
        data[175]=14;
        data[174]=14;
        data[173]=15;
        data[172]=15;
        data[171]=15;
        data[170]=16;
        data[169]=16;
        data[168]=17;
        data[167]=17;
        data[166]=17;
        data[165]=18;
        data[164]=18;
        data[163]=19;
        data[162]=19;
        data[161]=19;
        data[160]=20;
        data[159]=20;
        data[158]=21;
        data[157]=21;
        data[156]=22;
        data[155]=22;
        data[154]=23;
        data[153]=23;
        data[152]=24;
        data[151]=24;
        data[150]=24;
        data[149]=25;
        data[148]=25;
        data[147]=26;
        data[146]=26;
        data[145]=27;
        data[144]=27;
        data[143]=28;
        data[142]=28;
        data[141]=29;
        data[140]=29;
        data[139]=30;
        data[138]=30;
        data[137]=31;
        data[136]=31;
        data[135]=32;
        data[134]=33;
        data[133]=33;
        data[132]=34;
        data[131]=34;
        data[130]=35;
        data[129]=35;
        data[128]=36;
        data[127]=36;
        data[126]=37;
        data[125]=37;
        data[124]=38;
        data[123]=39;
        data[122]=39;
        data[121]=40;
        data[120]=40;
        data[119]=41;
        data[118]=42;
        data[117]=42;
        data[116]=43;
        data[115]=43;
        data[114]=44;
        data[113]=45;
        data[112]=45;
        data[111]=46;
        data[110]=46;
        data[109]=47;
        data[108]=48;
        data[107]=48;
        data[106]=49;
        data[105]=50;
        data[104]=50;
        data[103]=51;
        data[102]=51;
        data[101]=52;
        data[100]=53;
        data[99]=53;
        data[98]=54;
        data[97]=55;
        data[96]=55;
        data[95]=56;
        data[94]=57;
        data[93]=57;
        data[92]=58;
        data[91]=59;
        data[90]=59;
        data[89]=60;
        data[88]=61;
        data[87]=61;
        data[86]=62;
        data[85]=63;
        data[84]=64;
        data[83]=64;
        data[82]=65;
        data[81]=66;
        data[80]=66;
        data[79]=67;
        data[78]=68;
        data[77]=68;
        data[76]=69;
        data[75]=70;
        data[74]=71;
        data[73]=71;
        data[72]=72;
        data[71]=73;
        data[70]=74;
        data[69]=74;
        data[68]=75;
        data[67]=76;
        data[66]=76;
        data[65]=77;
        data[64]=78;
        data[63]=79;
        data[62]=79;
        data[61]=80;
        data[60]=81;
        data[59]=82;
        data[58]=82;
        data[57]=83;
        data[56]=84;
        data[55]=85;
        data[54]=85;
        data[53]=86;
        data[52]=87;
        data[51]=88;
        data[50]=88;
        data[49]=89;
        data[48]=90;
        data[47]=91;
        data[46]=92;
        data[45]=92;
        data[44]=93;
        data[43]=94;
        data[42]=95;
        data[41]=95;
        data[40]=96;
        data[39]=97;
        data[38]=98;
        data[37]=99;
        data[36]=99;
        data[35]=100;
        data[34]=101;
        data[33]=102;
        data[32]=102;
        data[31]=103;
        data[30]=104;
        data[29]=105;
        data[28]=106;
        data[27]=106;
        data[26]=107;
        data[25]=108;
        data[24]=109;
        data[23]=110;
        data[22]=110;
        data[21]=111;
        data[20]=112;
        data[19]=113;
        data[18]=114;
        data[17]=114;
        data[16]=115;
        data[15]=116;
        data[14]=117;
        data[13]=118;
        data[12]=118;
        data[11]=119;
        data[10]=120;
        data[9]=121;
        data[8]=122;
        data[7]=122;
        data[6]=123;
        data[5]=124;
        data[4]=125;
        data[3]=126;
        data[2]=126;
        data[1]=127;
        data[0]=128;

    end
    always @(posedge clk) begin
        
         otp<=data[{choose,count}];
        count<=(count+1'b1)%mod;
    end
    always @(posedge clk) begin
        if(count==999) cout<=1;
        else cout<=0;
    end
endmodule