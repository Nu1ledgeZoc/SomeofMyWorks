module rom2 (
    clk,
    otp
);
    input clk;
    output reg[7:0]otp;
    reg [7:0] data[999:0];
    reg [9:0] count;
    reg [9:0] mod;
    initial begin
         count=0;
        mod=1000;
        data[999]=255;
        data[998]=255;
        data[997]=255;
        data[996]=255;
        data[995]=255;
        data[994]=255;
        data[993]=255;
        data[992]=255;
        data[991]=255;
        data[990]=255;
        data[989]=255;
        data[988]=255;
        data[987]=255;
        data[986]=255;
        data[985]=255;
        data[984]=255;
        data[983]=255;
        data[982]=255;
        data[981]=255;
        data[980]=255;
        data[979]=255;
        data[978]=255;
        data[977]=255;
        data[976]=255;
        data[975]=255;
        data[974]=255;
        data[973]=255;
        data[972]=255;
        data[971]=255;
        data[970]=255;
        data[969]=255;
        data[968]=255;
        data[967]=255;
        data[966]=255;
        data[965]=255;
        data[964]=255;
        data[963]=255;
        data[962]=255;
        data[961]=255;
        data[960]=255;
        data[959]=255;
        data[958]=255;
        data[957]=255;
        data[956]=255;
        data[955]=255;
        data[954]=255;
        data[953]=255;
        data[952]=255;
        data[951]=255;
        data[950]=255;
        data[949]=255;
        data[948]=255;
        data[947]=255;
        data[946]=255;
        data[945]=255;
        data[944]=255;
        data[943]=255;
        data[942]=255;
        data[941]=255;
        data[940]=255;
        data[939]=255;
        data[938]=255;
        data[937]=255;
        data[936]=255;
        data[935]=255;
        data[934]=255;
        data[933]=255;
        data[932]=255;
        data[931]=255;
        data[930]=255;
        data[929]=255;
        data[928]=255;
        data[927]=255;
        data[926]=255;
        data[925]=255;
        data[924]=255;
        data[923]=255;
        data[922]=255;
        data[921]=255;
        data[920]=255;
        data[919]=255;
        data[918]=255;
        data[917]=255;
        data[916]=255;
        data[915]=255;
        data[914]=255;
        data[913]=255;
        data[912]=255;
        data[911]=255;
        data[910]=255;
        data[909]=255;
        data[908]=255;
        data[907]=255;
        data[906]=255;
        data[905]=255;
        data[904]=255;
        data[903]=255;
        data[902]=255;
        data[901]=255;
        data[900]=255;
        data[899]=255;
        data[898]=255;
        data[897]=255;
        data[896]=255;
        data[895]=255;
        data[894]=255;
        data[893]=255;
        data[892]=255;
        data[891]=255;
        data[890]=255;
        data[889]=255;
        data[888]=255;
        data[887]=255;
        data[886]=255;
        data[885]=255;
        data[884]=255;
        data[883]=255;
        data[882]=255;
        data[881]=255;
        data[880]=255;
        data[879]=255;
        data[878]=255;
        data[877]=255;
        data[876]=255;
        data[875]=255;
        data[874]=255;
        data[873]=255;
        data[872]=255;
        data[871]=255;
        data[870]=255;
        data[869]=255;
        data[868]=255;
        data[867]=255;
        data[866]=255;
        data[865]=255;
        data[864]=255;
        data[863]=255;
        data[862]=255;
        data[861]=255;
        data[860]=255;
        data[859]=255;
        data[858]=255;
        data[857]=255;
        data[856]=255;
        data[855]=255;
        data[854]=255;
        data[853]=255;
        data[852]=255;
        data[851]=255;
        data[850]=255;
        data[849]=255;
        data[848]=255;
        data[847]=255;
        data[846]=255;
        data[845]=255;
        data[844]=255;
        data[843]=255;
        data[842]=255;
        data[841]=255;
        data[840]=255;
        data[839]=255;
        data[838]=255;
        data[837]=255;
        data[836]=255;
        data[835]=255;
        data[834]=255;
        data[833]=255;
        data[832]=255;
        data[831]=255;
        data[830]=255;
        data[829]=255;
        data[828]=255;
        data[827]=255;
        data[826]=255;
        data[825]=255;
        data[824]=255;
        data[823]=255;
        data[822]=255;
        data[821]=255;
        data[820]=255;
        data[819]=255;
        data[818]=255;
        data[817]=255;
        data[816]=255;
        data[815]=255;
        data[814]=255;
        data[813]=255;
        data[812]=255;
        data[811]=255;
        data[810]=255;
        data[809]=255;
        data[808]=255;
        data[807]=255;
        data[806]=255;
        data[805]=255;
        data[804]=255;
        data[803]=255;
        data[802]=255;
        data[801]=255;
        data[800]=255;
        data[799]=255;
        data[798]=255;
        data[797]=255;
        data[796]=255;
        data[795]=255;
        data[794]=255;
        data[793]=255;
        data[792]=255;
        data[791]=255;
        data[790]=255;
        data[789]=255;
        data[788]=255;
        data[787]=255;
        data[786]=255;
        data[785]=255;
        data[784]=255;
        data[783]=255;
        data[782]=255;
        data[781]=255;
        data[780]=255;
        data[779]=255;
        data[778]=255;
        data[777]=255;
        data[776]=255;
        data[775]=255;
        data[774]=255;
        data[773]=255;
        data[772]=255;
        data[771]=255;
        data[770]=255;
        data[769]=255;
        data[768]=255;
        data[767]=255;
        data[766]=255;
        data[765]=255;
        data[764]=255;
        data[763]=255;
        data[762]=255;
        data[761]=255;
        data[760]=255;
        data[759]=255;
        data[758]=255;
        data[757]=255;
        data[756]=255;
        data[755]=255;
        data[754]=255;
        data[753]=255;
        data[752]=255;
        data[751]=255;
        data[750]=255;
        data[749]=255;
        data[748]=255;
        data[747]=255;
        data[746]=255;
        data[745]=255;
        data[744]=255;
        data[743]=255;
        data[742]=255;
        data[741]=255;
        data[740]=255;
        data[739]=255;
        data[738]=255;
        data[737]=255;
        data[736]=255;
        data[735]=255;
        data[734]=255;
        data[733]=255;
        data[732]=255;
        data[731]=255;
        data[730]=255;
        data[729]=255;
        data[728]=255;
        data[727]=255;
        data[726]=255;
        data[725]=255;
        data[724]=255;
        data[723]=255;
        data[722]=255;
        data[721]=255;
        data[720]=255;
        data[719]=255;
        data[718]=255;
        data[717]=255;
        data[716]=255;
        data[715]=255;
        data[714]=255;
        data[713]=255;
        data[712]=255;
        data[711]=255;
        data[710]=255;
        data[709]=255;
        data[708]=255;
        data[707]=255;
        data[706]=255;
        data[705]=255;
        data[704]=255;
        data[703]=255;
        data[702]=255;
        data[701]=255;
        data[700]=255;
        data[699]=255;
        data[698]=255;
        data[697]=255;
        data[696]=255;
        data[695]=255;
        data[694]=255;
        data[693]=255;
        data[692]=255;
        data[691]=255;
        data[690]=255;
        data[689]=255;
        data[688]=255;
        data[687]=255;
        data[686]=255;
        data[685]=255;
        data[684]=255;
        data[683]=255;
        data[682]=255;
        data[681]=255;
        data[680]=255;
        data[679]=255;
        data[678]=255;
        data[677]=255;
        data[676]=255;
        data[675]=255;
        data[674]=255;
        data[673]=255;
        data[672]=255;
        data[671]=255;
        data[670]=255;
        data[669]=255;
        data[668]=255;
        data[667]=255;
        data[666]=255;
        data[665]=255;
        data[664]=255;
        data[663]=255;
        data[662]=255;
        data[661]=255;
        data[660]=255;
        data[659]=255;
        data[658]=255;
        data[657]=255;
        data[656]=255;
        data[655]=255;
        data[654]=255;
        data[653]=255;
        data[652]=255;
        data[651]=255;
        data[650]=255;
        data[649]=255;
        data[648]=255;
        data[647]=255;
        data[646]=255;
        data[645]=255;
        data[644]=255;
        data[643]=255;
        data[642]=255;
        data[641]=255;
        data[640]=255;
        data[639]=255;
        data[638]=255;
        data[637]=255;
        data[636]=255;
        data[635]=255;
        data[634]=255;
        data[633]=255;
        data[632]=255;
        data[631]=255;
        data[630]=255;
        data[629]=255;
        data[628]=255;
        data[627]=255;
        data[626]=255;
        data[625]=255;
        data[624]=255;
        data[623]=255;
        data[622]=255;
        data[621]=255;
        data[620]=255;
        data[619]=255;
        data[618]=255;
        data[617]=255;
        data[616]=255;
        data[615]=255;
        data[614]=255;
        data[613]=255;
        data[612]=255;
        data[611]=255;
        data[610]=255;
        data[609]=255;
        data[608]=255;
        data[607]=255;
        data[606]=255;
        data[605]=255;
        data[604]=255;
        data[603]=255;
        data[602]=255;
        data[601]=255;
        data[600]=255;
        data[599]=255;
        data[598]=255;
        data[597]=255;
        data[596]=255;
        data[595]=255;
        data[594]=255;
        data[593]=255;
        data[592]=255;
        data[591]=255;
        data[590]=255;
        data[589]=255;
        data[588]=255;
        data[587]=255;
        data[586]=255;
        data[585]=255;
        data[584]=255;
        data[583]=255;
        data[582]=255;
        data[581]=255;
        data[580]=255;
        data[579]=255;
        data[578]=255;
        data[577]=255;
        data[576]=255;
        data[575]=255;
        data[574]=255;
        data[573]=255;
        data[572]=255;
        data[571]=255;
        data[570]=255;
        data[569]=255;
        data[568]=255;
        data[567]=255;
        data[566]=255;
        data[565]=255;
        data[564]=255;
        data[563]=255;
        data[562]=255;
        data[561]=255;
        data[560]=255;
        data[559]=255;
        data[558]=255;
        data[557]=255;
        data[556]=255;
        data[555]=255;
        data[554]=255;
        data[553]=255;
        data[552]=255;
        data[551]=255;
        data[550]=255;
        data[549]=255;
        data[548]=255;
        data[547]=255;
        data[546]=255;
        data[545]=255;
        data[544]=255;
        data[543]=255;
        data[542]=255;
        data[541]=255;
        data[540]=255;
        data[539]=255;
        data[538]=255;
        data[537]=255;
        data[536]=255;
        data[535]=255;
        data[534]=255;
        data[533]=255;
        data[532]=255;
        data[531]=255;
        data[530]=255;
        data[529]=255;
        data[528]=255;
        data[527]=255;
        data[526]=255;
        data[525]=255;
        data[524]=255;
        data[523]=255;
        data[522]=255;
        data[521]=255;
        data[520]=255;
        data[519]=255;
        data[518]=255;
        data[517]=255;
        data[516]=255;
        data[515]=255;
        data[514]=255;
        data[513]=255;
        data[512]=255;
        data[511]=255;
        data[510]=255;
        data[509]=255;
        data[508]=255;
        data[507]=255;
        data[506]=255;
        data[505]=255;
        data[504]=255;
        data[503]=255;
        data[502]=255;
        data[501]=255;
        data[500]=255;
        data[499]=0;
        data[498]=0;
        data[497]=0;
        data[496]=0;
        data[495]=0;
        data[494]=0;
        data[493]=0;
        data[492]=0;
        data[491]=0;
        data[490]=0;
        data[489]=0;
        data[488]=0;
        data[487]=0;
        data[486]=0;
        data[485]=0;
        data[484]=0;
        data[483]=0;
        data[482]=0;
        data[481]=0;
        data[480]=0;
        data[479]=0;
        data[478]=0;
        data[477]=0;
        data[476]=0;
        data[475]=0;
        data[474]=0;
        data[473]=0;
        data[472]=0;
        data[471]=0;
        data[470]=0;
        data[469]=0;
        data[468]=0;
        data[467]=0;
        data[466]=0;
        data[465]=0;
        data[464]=0;
        data[463]=0;
        data[462]=0;
        data[461]=0;
        data[460]=0;
        data[459]=0;
        data[458]=0;
        data[457]=0;
        data[456]=0;
        data[455]=0;
        data[454]=0;
        data[453]=0;
        data[452]=0;
        data[451]=0;
        data[450]=0;
        data[449]=0;
        data[448]=0;
        data[447]=0;
        data[446]=0;
        data[445]=0;
        data[444]=0;
        data[443]=0;
        data[442]=0;
        data[441]=0;
        data[440]=0;
        data[439]=0;
        data[438]=0;
        data[437]=0;
        data[436]=0;
        data[435]=0;
        data[434]=0;
        data[433]=0;
        data[432]=0;
        data[431]=0;
        data[430]=0;
        data[429]=0;
        data[428]=0;
        data[427]=0;
        data[426]=0;
        data[425]=0;
        data[424]=0;
        data[423]=0;
        data[422]=0;
        data[421]=0;
        data[420]=0;
        data[419]=0;
        data[418]=0;
        data[417]=0;
        data[416]=0;
        data[415]=0;
        data[414]=0;
        data[413]=0;
        data[412]=0;
        data[411]=0;
        data[410]=0;
        data[409]=0;
        data[408]=0;
        data[407]=0;
        data[406]=0;
        data[405]=0;
        data[404]=0;
        data[403]=0;
        data[402]=0;
        data[401]=0;
        data[400]=0;
        data[399]=0;
        data[398]=0;
        data[397]=0;
        data[396]=0;
        data[395]=0;
        data[394]=0;
        data[393]=0;
        data[392]=0;
        data[391]=0;
        data[390]=0;
        data[389]=0;
        data[388]=0;
        data[387]=0;
        data[386]=0;
        data[385]=0;
        data[384]=0;
        data[383]=0;
        data[382]=0;
        data[381]=0;
        data[380]=0;
        data[379]=0;
        data[378]=0;
        data[377]=0;
        data[376]=0;
        data[375]=0;
        data[374]=0;
        data[373]=0;
        data[372]=0;
        data[371]=0;
        data[370]=0;
        data[369]=0;
        data[368]=0;
        data[367]=0;
        data[366]=0;
        data[365]=0;
        data[364]=0;
        data[363]=0;
        data[362]=0;
        data[361]=0;
        data[360]=0;
        data[359]=0;
        data[358]=0;
        data[357]=0;
        data[356]=0;
        data[355]=0;
        data[354]=0;
        data[353]=0;
        data[352]=0;
        data[351]=0;
        data[350]=0;
        data[349]=0;
        data[348]=0;
        data[347]=0;
        data[346]=0;
        data[345]=0;
        data[344]=0;
        data[343]=0;
        data[342]=0;
        data[341]=0;
        data[340]=0;
        data[339]=0;
        data[338]=0;
        data[337]=0;
        data[336]=0;
        data[335]=0;
        data[334]=0;
        data[333]=0;
        data[332]=0;
        data[331]=0;
        data[330]=0;
        data[329]=0;
        data[328]=0;
        data[327]=0;
        data[326]=0;
        data[325]=0;
        data[324]=0;
        data[323]=0;
        data[322]=0;
        data[321]=0;
        data[320]=0;
        data[319]=0;
        data[318]=0;
        data[317]=0;
        data[316]=0;
        data[315]=0;
        data[314]=0;
        data[313]=0;
        data[312]=0;
        data[311]=0;
        data[310]=0;
        data[309]=0;
        data[308]=0;
        data[307]=0;
        data[306]=0;
        data[305]=0;
        data[304]=0;
        data[303]=0;
        data[302]=0;
        data[301]=0;
        data[300]=0;
        data[299]=0;
        data[298]=0;
        data[297]=0;
        data[296]=0;
        data[295]=0;
        data[294]=0;
        data[293]=0;
        data[292]=0;
        data[291]=0;
        data[290]=0;
        data[289]=0;
        data[288]=0;
        data[287]=0;
        data[286]=0;
        data[285]=0;
        data[284]=0;
        data[283]=0;
        data[282]=0;
        data[281]=0;
        data[280]=0;
        data[279]=0;
        data[278]=0;
        data[277]=0;
        data[276]=0;
        data[275]=0;
        data[274]=0;
        data[273]=0;
        data[272]=0;
        data[271]=0;
        data[270]=0;
        data[269]=0;
        data[268]=0;
        data[267]=0;
        data[266]=0;
        data[265]=0;
        data[264]=0;
        data[263]=0;
        data[262]=0;
        data[261]=0;
        data[260]=0;
        data[259]=0;
        data[258]=0;
        data[257]=0;
        data[256]=0;
        data[255]=0;
        data[254]=0;
        data[253]=0;
        data[252]=0;
        data[251]=0;
        data[250]=0;
        data[249]=0;
        data[248]=0;
        data[247]=0;
        data[246]=0;
        data[245]=0;
        data[244]=0;
        data[243]=0;
        data[242]=0;
        data[241]=0;
        data[240]=0;
        data[239]=0;
        data[238]=0;
        data[237]=0;
        data[236]=0;
        data[235]=0;
        data[234]=0;
        data[233]=0;
        data[232]=0;
        data[231]=0;
        data[230]=0;
        data[229]=0;
        data[228]=0;
        data[227]=0;
        data[226]=0;
        data[225]=0;
        data[224]=0;
        data[223]=0;
        data[222]=0;
        data[221]=0;
        data[220]=0;
        data[219]=0;
        data[218]=0;
        data[217]=0;
        data[216]=0;
        data[215]=0;
        data[214]=0;
        data[213]=0;
        data[212]=0;
        data[211]=0;
        data[210]=0;
        data[209]=0;
        data[208]=0;
        data[207]=0;
        data[206]=0;
        data[205]=0;
        data[204]=0;
        data[203]=0;
        data[202]=0;
        data[201]=0;
        data[200]=0;
        data[199]=0;
        data[198]=0;
        data[197]=0;
        data[196]=0;
        data[195]=0;
        data[194]=0;
        data[193]=0;
        data[192]=0;
        data[191]=0;
        data[190]=0;
        data[189]=0;
        data[188]=0;
        data[187]=0;
        data[186]=0;
        data[185]=0;
        data[184]=0;
        data[183]=0;
        data[182]=0;
        data[181]=0;
        data[180]=0;
        data[179]=0;
        data[178]=0;
        data[177]=0;
        data[176]=0;
        data[175]=0;
        data[174]=0;
        data[173]=0;
        data[172]=0;
        data[171]=0;
        data[170]=0;
        data[169]=0;
        data[168]=0;
        data[167]=0;
        data[166]=0;
        data[165]=0;
        data[164]=0;
        data[163]=0;
        data[162]=0;
        data[161]=0;
        data[160]=0;
        data[159]=0;
        data[158]=0;
        data[157]=0;
        data[156]=0;
        data[155]=0;
        data[154]=0;
        data[153]=0;
        data[152]=0;
        data[151]=0;
        data[150]=0;
        data[149]=0;
        data[148]=0;
        data[147]=0;
        data[146]=0;
        data[145]=0;
        data[144]=0;
        data[143]=0;
        data[142]=0;
        data[141]=0;
        data[140]=0;
        data[139]=0;
        data[138]=0;
        data[137]=0;
        data[136]=0;
        data[135]=0;
        data[134]=0;
        data[133]=0;
        data[132]=0;
        data[131]=0;
        data[130]=0;
        data[129]=0;
        data[128]=0;
        data[127]=0;
        data[126]=0;
        data[125]=0;
        data[124]=0;
        data[123]=0;
        data[122]=0;
        data[121]=0;
        data[120]=0;
        data[119]=0;
        data[118]=0;
        data[117]=0;
        data[116]=0;
        data[115]=0;
        data[114]=0;
        data[113]=0;
        data[112]=0;
        data[111]=0;
        data[110]=0;
        data[109]=0;
        data[108]=0;
        data[107]=0;
        data[106]=0;
        data[105]=0;
        data[104]=0;
        data[103]=0;
        data[102]=0;
        data[101]=0;
        data[100]=0;
        data[99]=0;
        data[98]=0;
        data[97]=0;
        data[96]=0;
        data[95]=0;
        data[94]=0;
        data[93]=0;
        data[92]=0;
        data[91]=0;
        data[90]=0;
        data[89]=0;
        data[88]=0;
        data[87]=0;
        data[86]=0;
        data[85]=0;
        data[84]=0;
        data[83]=0;
        data[82]=0;
        data[81]=0;
        data[80]=0;
        data[79]=0;
        data[78]=0;
        data[77]=0;
        data[76]=0;
        data[75]=0;
        data[74]=0;
        data[73]=0;
        data[72]=0;
        data[71]=0;
        data[70]=0;
        data[69]=0;
        data[68]=0;
        data[67]=0;
        data[66]=0;
        data[65]=0;
        data[64]=0;
        data[63]=0;
        data[62]=0;
        data[61]=0;
        data[60]=0;
        data[59]=0;
        data[58]=0;
        data[57]=0;
        data[56]=0;
        data[55]=0;
        data[54]=0;
        data[53]=0;
        data[52]=0;
        data[51]=0;
        data[50]=0;
        data[49]=0;
        data[48]=0;
        data[47]=0;
        data[46]=0;
        data[45]=0;
        data[44]=0;
        data[43]=0;
        data[42]=0;
        data[41]=0;
        data[40]=0;
        data[39]=0;
        data[38]=0;
        data[37]=0;
        data[36]=0;
        data[35]=0;
        data[34]=0;
        data[33]=0;
        data[32]=0;
        data[31]=0;
        data[30]=0;
        data[29]=0;
        data[28]=0;
        data[27]=0;
        data[26]=0;
        data[25]=0;
        data[24]=0;
        data[23]=0;
        data[22]=0;
        data[21]=0;
        data[20]=0;
        data[19]=0;
        data[18]=0;
        data[17]=0;
        data[16]=0;
        data[15]=0;
        data[14]=0;
        data[13]=0;
        data[12]=0;
        data[11]=0;
        data[10]=0;
        data[9]=0;
        data[8]=0;
        data[7]=0;
        data[6]=0;
        data[5]=0;
        data[4]=0;
        data[3]=0;
        data[2]=0;
        data[1]=0;
        data[0]=0;

    end
     always @(posedge clk) begin
        otp<=data[count];
        count<=(count+1'b1)%mod;
    end
endmodule