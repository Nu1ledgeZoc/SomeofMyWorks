module rom4 (
    clk,
    otp
);
    input clk;
    output reg[7:0]otp;
    reg [7:0] data[999:0];
    reg [9:0] count;
    reg [9:0] mod;
    initial begin
         count=0;
        mod=1000;
        data[999]=0;
        data[998]=3;
        data[997]=5;
        data[996]=8;
        data[995]=10;
        data[994]=13;
        data[993]=15;
        data[992]=18;
        data[991]=20;
        data[990]=23;
        data[989]=25;
        data[988]=28;
        data[987]=31;
        data[986]=33;
        data[985]=36;
        data[984]=38;
        data[983]=41;
        data[982]=43;
        data[981]=46;
        data[980]=48;
        data[979]=51;
        data[978]=54;
        data[977]=56;
        data[976]=59;
        data[975]=61;
        data[974]=64;
        data[973]=66;
        data[972]=69;
        data[971]=71;
        data[970]=74;
        data[969]=77;
        data[968]=79;
        data[967]=82;
        data[966]=84;
        data[965]=87;
        data[964]=89;
        data[963]=92;
        data[962]=94;
        data[961]=97;
        data[960]=99;
        data[959]=102;
        data[958]=105;
        data[957]=107;
        data[956]=110;
        data[955]=112;
        data[954]=115;
        data[953]=117;
        data[952]=120;
        data[951]=122;
        data[950]=125;
        data[949]=127;
        data[948]=130;
        data[947]=133;
        data[946]=135;
        data[945]=138;
        data[944]=140;
        data[943]=143;
        data[942]=145;
        data[941]=148;
        data[940]=150;
        data[939]=153;
        data[938]=156;
        data[937]=158;
        data[936]=161;
        data[935]=163;
        data[934]=166;
        data[933]=168;
        data[932]=171;
        data[931]=173;
        data[930]=176;
        data[929]=179;
        data[928]=181;
        data[927]=184;
        data[926]=186;
        data[925]=189;
        data[924]=191;
        data[923]=194;
        data[922]=196;
        data[921]=199;
        data[920]=201;
        data[919]=204;
        data[918]=207;
        data[917]=209;
        data[916]=212;
        data[915]=214;
        data[914]=217;
        data[913]=219;
        data[912]=222;
        data[911]=224;
        data[910]=227;
        data[909]=229;
        data[908]=232;
        data[907]=235;
        data[906]=237;
        data[905]=240;
        data[904]=242;
        data[903]=245;
        data[902]=247;
        data[901]=250;
        data[900]=252;
        data[899]=255;
        data[898]=254;
        data[897]=254;
        data[896]=254;
        data[895]=254;
        data[894]=253;
        data[893]=253;
        data[892]=253;
        data[891]=252;
        data[890]=252;
        data[889]=252;
        data[888]=252;
        data[887]=251;
        data[886]=251;
        data[885]=251;
        data[884]=250;
        data[883]=250;
        data[882]=250;
        data[881]=250;
        data[880]=249;
        data[879]=249;
        data[878]=249;
        data[877]=248;
        data[876]=248;
        data[875]=248;
        data[874]=248;
        data[873]=247;
        data[872]=247;
        data[871]=247;
        data[870]=247;
        data[869]=246;
        data[868]=246;
        data[867]=246;
        data[866]=245;
        data[865]=245;
        data[864]=245;
        data[863]=245;
        data[862]=244;
        data[861]=244;
        data[860]=244;
        data[859]=243;
        data[858]=243;
        data[857]=243;
        data[856]=243;
        data[855]=242;
        data[854]=242;
        data[853]=242;
        data[852]=241;
        data[851]=241;
        data[850]=241;
        data[849]=241;
        data[848]=240;
        data[847]=240;
        data[846]=240;
        data[845]=239;
        data[844]=239;
        data[843]=239;
        data[842]=239;
        data[841]=238;
        data[840]=238;
        data[839]=238;
        data[838]=237;
        data[837]=237;
        data[836]=237;
        data[835]=237;
        data[834]=236;
        data[833]=236;
        data[832]=236;
        data[831]=235;
        data[830]=235;
        data[829]=235;
        data[828]=235;
        data[827]=234;
        data[826]=234;
        data[825]=234;
        data[824]=233;
        data[823]=233;
        data[822]=233;
        data[821]=233;
        data[820]=232;
        data[819]=232;
        data[818]=232;
        data[817]=231;
        data[816]=231;
        data[815]=231;
        data[814]=231;
        data[813]=230;
        data[812]=230;
        data[811]=230;
        data[810]=229;
        data[809]=229;
        data[808]=229;
        data[807]=229;
        data[806]=228;
        data[805]=228;
        data[804]=228;
        data[803]=228;
        data[802]=227;
        data[801]=227;
        data[800]=227;
        data[799]=226;
        data[798]=226;
        data[797]=226;
        data[796]=226;
        data[795]=225;
        data[794]=225;
        data[793]=225;
        data[792]=224;
        data[791]=224;
        data[790]=224;
        data[789]=224;
        data[788]=223;
        data[787]=223;
        data[786]=223;
        data[785]=222;
        data[784]=222;
        data[783]=222;
        data[782]=222;
        data[781]=221;
        data[780]=221;
        data[779]=221;
        data[778]=220;
        data[777]=220;
        data[776]=220;
        data[775]=220;
        data[774]=219;
        data[773]=219;
        data[772]=219;
        data[771]=218;
        data[770]=218;
        data[769]=218;
        data[768]=218;
        data[767]=217;
        data[766]=217;
        data[765]=217;
        data[764]=216;
        data[763]=216;
        data[762]=216;
        data[761]=216;
        data[760]=215;
        data[759]=215;
        data[758]=215;
        data[757]=214;
        data[756]=214;
        data[755]=214;
        data[754]=214;
        data[753]=213;
        data[752]=213;
        data[751]=213;
        data[750]=213;
        data[749]=212;
        data[748]=212;
        data[747]=212;
        data[746]=211;
        data[745]=211;
        data[744]=211;
        data[743]=211;
        data[742]=210;
        data[741]=210;
        data[740]=210;
        data[739]=209;
        data[738]=209;
        data[737]=209;
        data[736]=209;
        data[735]=208;
        data[734]=208;
        data[733]=208;
        data[732]=207;
        data[731]=207;
        data[730]=207;
        data[729]=207;
        data[728]=206;
        data[727]=206;
        data[726]=206;
        data[725]=205;
        data[724]=205;
        data[723]=205;
        data[722]=205;
        data[721]=204;
        data[720]=204;
        data[719]=204;
        data[718]=203;
        data[717]=203;
        data[716]=203;
        data[715]=203;
        data[714]=202;
        data[713]=202;
        data[712]=202;
        data[711]=201;
        data[710]=201;
        data[709]=201;
        data[708]=201;
        data[707]=200;
        data[706]=200;
        data[705]=200;
        data[704]=199;
        data[703]=199;
        data[702]=199;
        data[701]=199;
        data[700]=198;
        data[699]=198;
        data[698]=198;
        data[697]=197;
        data[696]=197;
        data[695]=197;
        data[694]=197;
        data[693]=196;
        data[692]=196;
        data[691]=196;
        data[690]=195;
        data[689]=195;
        data[688]=195;
        data[687]=195;
        data[686]=194;
        data[685]=194;
        data[684]=194;
        data[683]=194;
        data[682]=193;
        data[681]=193;
        data[680]=193;
        data[679]=192;
        data[678]=192;
        data[677]=192;
        data[676]=192;
        data[675]=191;
        data[674]=191;
        data[673]=191;
        data[672]=190;
        data[671]=190;
        data[670]=190;
        data[669]=190;
        data[668]=189;
        data[667]=189;
        data[666]=189;
        data[665]=188;
        data[664]=188;
        data[663]=188;
        data[662]=188;
        data[661]=187;
        data[660]=187;
        data[659]=187;
        data[658]=186;
        data[657]=186;
        data[656]=186;
        data[655]=186;
        data[654]=185;
        data[653]=185;
        data[652]=185;
        data[651]=184;
        data[650]=184;
        data[649]=184;
        data[648]=184;
        data[647]=183;
        data[646]=183;
        data[645]=183;
        data[644]=182;
        data[643]=182;
        data[642]=182;
        data[641]=182;
        data[640]=181;
        data[639]=181;
        data[638]=181;
        data[637]=180;
        data[636]=180;
        data[635]=180;
        data[634]=180;
        data[633]=179;
        data[632]=179;
        data[631]=179;
        data[630]=178;
        data[629]=178;
        data[628]=178;
        data[627]=178;
        data[626]=177;
        data[625]=177;
        data[624]=177;
        data[623]=177;
        data[622]=176;
        data[621]=176;
        data[620]=176;
        data[619]=175;
        data[618]=175;
        data[617]=175;
        data[616]=175;
        data[615]=174;
        data[614]=174;
        data[613]=174;
        data[612]=173;
        data[611]=173;
        data[610]=173;
        data[609]=173;
        data[608]=172;
        data[607]=172;
        data[606]=172;
        data[605]=171;
        data[604]=171;
        data[603]=171;
        data[602]=171;
        data[601]=170;
        data[600]=170;
        data[599]=170;
        data[598]=169;
        data[597]=169;
        data[596]=169;
        data[595]=169;
        data[594]=168;
        data[593]=168;
        data[592]=168;
        data[591]=167;
        data[590]=167;
        data[589]=167;
        data[588]=167;
        data[587]=166;
        data[586]=166;
        data[585]=166;
        data[584]=165;
        data[583]=165;
        data[582]=165;
        data[581]=165;
        data[580]=164;
        data[579]=164;
        data[578]=164;
        data[577]=163;
        data[576]=163;
        data[575]=163;
        data[574]=163;
        data[573]=162;
        data[572]=162;
        data[571]=162;
        data[570]=162;
        data[569]=161;
        data[568]=161;
        data[567]=161;
        data[566]=160;
        data[565]=160;
        data[564]=160;
        data[563]=160;
        data[562]=159;
        data[561]=159;
        data[560]=159;
        data[559]=158;
        data[558]=158;
        data[557]=158;
        data[556]=158;
        data[555]=157;
        data[554]=157;
        data[553]=157;
        data[552]=156;
        data[551]=156;
        data[550]=156;
        data[549]=156;
        data[548]=155;
        data[547]=155;
        data[546]=155;
        data[545]=154;
        data[544]=154;
        data[543]=154;
        data[542]=154;
        data[541]=153;
        data[540]=153;
        data[539]=153;
        data[538]=152;
        data[537]=152;
        data[536]=152;
        data[535]=152;
        data[534]=151;
        data[533]=151;
        data[532]=151;
        data[531]=150;
        data[530]=150;
        data[529]=150;
        data[528]=150;
        data[527]=149;
        data[526]=149;
        data[525]=149;
        data[524]=148;
        data[523]=148;
        data[522]=148;
        data[521]=148;
        data[520]=147;
        data[519]=147;
        data[518]=147;
        data[517]=146;
        data[516]=146;
        data[515]=146;
        data[514]=146;
        data[513]=145;
        data[512]=145;
        data[511]=145;
        data[510]=144;
        data[509]=144;
        data[508]=144;
        data[507]=144;
        data[506]=143;
        data[505]=143;
        data[504]=143;
        data[503]=143;
        data[502]=142;
        data[501]=142;
        data[500]=142;
        data[499]=141;
        data[498]=141;
        data[497]=141;
        data[496]=141;
        data[495]=140;
        data[494]=140;
        data[493]=140;
        data[492]=139;
        data[491]=139;
        data[490]=139;
        data[489]=139;
        data[488]=138;
        data[487]=138;
        data[486]=138;
        data[485]=137;
        data[484]=137;
        data[483]=137;
        data[482]=137;
        data[481]=136;
        data[480]=136;
        data[479]=136;
        data[478]=135;
        data[477]=135;
        data[476]=135;
        data[475]=135;
        data[474]=134;
        data[473]=134;
        data[472]=134;
        data[471]=133;
        data[470]=133;
        data[469]=133;
        data[468]=133;
        data[467]=132;
        data[466]=132;
        data[465]=132;
        data[464]=131;
        data[463]=131;
        data[462]=131;
        data[461]=131;
        data[460]=130;
        data[459]=130;
        data[458]=130;
        data[457]=129;
        data[456]=129;
        data[455]=129;
        data[454]=129;
        data[453]=128;
        data[452]=128;
        data[451]=128;
        data[450]=128;
        data[449]=127;
        data[448]=127;
        data[447]=127;
        data[446]=126;
        data[445]=126;
        data[444]=126;
        data[443]=126;
        data[442]=125;
        data[441]=125;
        data[440]=125;
        data[439]=124;
        data[438]=124;
        data[437]=124;
        data[436]=124;
        data[435]=123;
        data[434]=123;
        data[433]=123;
        data[432]=122;
        data[431]=122;
        data[430]=122;
        data[429]=122;
        data[428]=121;
        data[427]=121;
        data[426]=121;
        data[425]=120;
        data[424]=120;
        data[423]=120;
        data[422]=120;
        data[421]=119;
        data[420]=119;
        data[419]=119;
        data[418]=118;
        data[417]=118;
        data[416]=118;
        data[415]=118;
        data[414]=117;
        data[413]=117;
        data[412]=117;
        data[411]=116;
        data[410]=116;
        data[409]=116;
        data[408]=116;
        data[407]=115;
        data[406]=115;
        data[405]=115;
        data[404]=114;
        data[403]=114;
        data[402]=114;
        data[401]=114;
        data[400]=113;
        data[399]=113;
        data[398]=113;
        data[397]=112;
        data[396]=112;
        data[395]=112;
        data[394]=112;
        data[393]=111;
        data[392]=111;
        data[391]=111;
        data[390]=110;
        data[389]=110;
        data[388]=110;
        data[387]=110;
        data[386]=109;
        data[385]=109;
        data[384]=109;
        data[383]=109;
        data[382]=108;
        data[381]=108;
        data[380]=108;
        data[379]=107;
        data[378]=107;
        data[377]=107;
        data[376]=107;
        data[375]=106;
        data[374]=106;
        data[373]=106;
        data[372]=105;
        data[371]=105;
        data[370]=105;
        data[369]=105;
        data[368]=104;
        data[367]=104;
        data[366]=104;
        data[365]=103;
        data[364]=103;
        data[363]=103;
        data[362]=103;
        data[361]=102;
        data[360]=102;
        data[359]=102;
        data[358]=101;
        data[357]=101;
        data[356]=101;
        data[355]=101;
        data[354]=100;
        data[353]=100;
        data[352]=100;
        data[351]=99;
        data[350]=99;
        data[349]=99;
        data[348]=99;
        data[347]=98;
        data[346]=98;
        data[345]=98;
        data[344]=97;
        data[343]=97;
        data[342]=97;
        data[341]=97;
        data[340]=96;
        data[339]=96;
        data[338]=96;
        data[337]=95;
        data[336]=95;
        data[335]=95;
        data[334]=95;
        data[333]=94;
        data[332]=94;
        data[331]=94;
        data[330]=94;
        data[329]=93;
        data[328]=93;
        data[327]=93;
        data[326]=92;
        data[325]=92;
        data[324]=92;
        data[323]=92;
        data[322]=91;
        data[321]=91;
        data[320]=91;
        data[319]=90;
        data[318]=90;
        data[317]=90;
        data[316]=90;
        data[315]=89;
        data[314]=89;
        data[313]=89;
        data[312]=88;
        data[311]=88;
        data[310]=88;
        data[309]=88;
        data[308]=87;
        data[307]=87;
        data[306]=87;
        data[305]=86;
        data[304]=86;
        data[303]=86;
        data[302]=86;
        data[301]=85;
        data[300]=85;
        data[299]=85;
        data[298]=84;
        data[297]=84;
        data[296]=84;
        data[295]=84;
        data[294]=83;
        data[293]=83;
        data[292]=83;
        data[291]=82;
        data[290]=82;
        data[289]=82;
        data[288]=82;
        data[287]=81;
        data[286]=81;
        data[285]=81;
        data[284]=80;
        data[283]=80;
        data[282]=80;
        data[281]=80;
        data[280]=79;
        data[279]=79;
        data[278]=79;
        data[277]=78;
        data[276]=78;
        data[275]=78;
        data[274]=78;
        data[273]=77;
        data[272]=77;
        data[271]=77;
        data[270]=77;
        data[269]=76;
        data[268]=76;
        data[267]=76;
        data[266]=75;
        data[265]=75;
        data[264]=75;
        data[263]=75;
        data[262]=74;
        data[261]=74;
        data[260]=74;
        data[259]=73;
        data[258]=73;
        data[257]=73;
        data[256]=73;
        data[255]=72;
        data[254]=72;
        data[253]=72;
        data[252]=71;
        data[251]=71;
        data[250]=71;
        data[249]=71;
        data[248]=70;
        data[247]=70;
        data[246]=70;
        data[245]=69;
        data[244]=69;
        data[243]=69;
        data[242]=69;
        data[241]=68;
        data[240]=68;
        data[239]=68;
        data[238]=67;
        data[237]=67;
        data[236]=67;
        data[235]=67;
        data[234]=66;
        data[233]=66;
        data[232]=66;
        data[231]=65;
        data[230]=65;
        data[229]=65;
        data[228]=65;
        data[227]=64;
        data[226]=64;
        data[225]=64;
        data[224]=63;
        data[223]=63;
        data[222]=63;
        data[221]=63;
        data[220]=62;
        data[219]=62;
        data[218]=62;
        data[217]=61;
        data[216]=61;
        data[215]=61;
        data[214]=61;
        data[213]=60;
        data[212]=60;
        data[211]=60;
        data[210]=59;
        data[209]=59;
        data[208]=59;
        data[207]=59;
        data[206]=58;
        data[205]=58;
        data[204]=58;
        data[203]=58;
        data[202]=57;
        data[201]=57;
        data[200]=57;
        data[199]=56;
        data[198]=56;
        data[197]=56;
        data[196]=56;
        data[195]=55;
        data[194]=55;
        data[193]=55;
        data[192]=54;
        data[191]=54;
        data[190]=54;
        data[189]=54;
        data[188]=53;
        data[187]=53;
        data[186]=53;
        data[185]=52;
        data[184]=52;
        data[183]=52;
        data[182]=52;
        data[181]=51;
        data[180]=51;
        data[179]=51;
        data[178]=50;
        data[177]=50;
        data[176]=50;
        data[175]=50;
        data[174]=49;
        data[173]=49;
        data[172]=49;
        data[171]=48;
        data[170]=48;
        data[169]=48;
        data[168]=48;
        data[167]=47;
        data[166]=47;
        data[165]=47;
        data[164]=46;
        data[163]=46;
        data[162]=46;
        data[161]=46;
        data[160]=45;
        data[159]=45;
        data[158]=45;
        data[157]=44;
        data[156]=44;
        data[155]=44;
        data[154]=44;
        data[153]=43;
        data[152]=43;
        data[151]=43;
        data[150]=43;
        data[149]=42;
        data[148]=42;
        data[147]=42;
        data[146]=41;
        data[145]=41;
        data[144]=41;
        data[143]=41;
        data[142]=40;
        data[141]=40;
        data[140]=40;
        data[139]=39;
        data[138]=39;
        data[137]=39;
        data[136]=39;
        data[135]=38;
        data[134]=38;
        data[133]=38;
        data[132]=37;
        data[131]=37;
        data[130]=37;
        data[129]=37;
        data[128]=36;
        data[127]=36;
        data[126]=36;
        data[125]=35;
        data[124]=35;
        data[123]=35;
        data[122]=35;
        data[121]=34;
        data[120]=34;
        data[119]=34;
        data[118]=33;
        data[117]=33;
        data[116]=33;
        data[115]=33;
        data[114]=32;
        data[113]=32;
        data[112]=32;
        data[111]=31;
        data[110]=31;
        data[109]=31;
        data[108]=31;
        data[107]=30;
        data[106]=30;
        data[105]=30;
        data[104]=29;
        data[103]=29;
        data[102]=29;
        data[101]=29;
        data[100]=28;
        data[99]=28;
        data[98]=28;
        data[97]=27;
        data[96]=27;
        data[95]=27;
        data[94]=27;
        data[93]=26;
        data[92]=26;
        data[91]=26;
        data[90]=25;
        data[89]=25;
        data[88]=25;
        data[87]=25;
        data[86]=24;
        data[85]=24;
        data[84]=24;
        data[83]=24;
        data[82]=23;
        data[81]=23;
        data[80]=23;
        data[79]=22;
        data[78]=22;
        data[77]=22;
        data[76]=22;
        data[75]=21;
        data[74]=21;
        data[73]=21;
        data[72]=20;
        data[71]=20;
        data[70]=20;
        data[69]=20;
        data[68]=19;
        data[67]=19;
        data[66]=19;
        data[65]=18;
        data[64]=18;
        data[63]=18;
        data[62]=18;
        data[61]=17;
        data[60]=17;
        data[59]=17;
        data[58]=16;
        data[57]=16;
        data[56]=16;
        data[55]=16;
        data[54]=15;
        data[53]=15;
        data[52]=15;
        data[51]=14;
        data[50]=14;
        data[49]=14;
        data[48]=14;
        data[47]=13;
        data[46]=13;
        data[45]=13;
        data[44]=12;
        data[43]=12;
        data[42]=12;
        data[41]=12;
        data[40]=11;
        data[39]=11;
        data[38]=11;
        data[37]=10;
        data[36]=10;
        data[35]=10;
        data[34]=10;
        data[33]=9;
        data[32]=9;
        data[31]=9;
        data[30]=9;
        data[29]=8;
        data[28]=8;
        data[27]=8;
        data[26]=7;
        data[25]=7;
        data[24]=7;
        data[23]=7;
        data[22]=6;
        data[21]=6;
        data[20]=6;
        data[19]=5;
        data[18]=5;
        data[17]=5;
        data[16]=5;
        data[15]=4;
        data[14]=4;
        data[13]=4;
        data[12]=3;
        data[11]=3;
        data[10]=3;
        data[9]=3;
        data[8]=2;
        data[7]=2;
        data[6]=2;
        data[5]=1;
        data[4]=1;
        data[3]=1;
        data[2]=1;
        data[1]=0;
        data[0]=0;

    end
     always @(posedge clk) begin
        otp<=data[count];
        count<=(count+1'b1)%mod;
    end
endmodule