module romtatal (
    clk,
    choose,
    cout,
    otp
);
    input clk;
    input [1:0] choose;
    output reg[7:0] otp;
    output reg cout;
    reg [7:0] data[4095:0];
    reg [9:0] count;
    reg [9:0] mod;
   
    initial begin
        cout=0;
         otp=0;
         count=0;
        mod=1000;
        data[4095]=0;
        data[4094]=0;
        data[4093]=0;
        data[4092]=0;
        data[4091]=0;
        data[4090]=0;
        data[4089]=0;
        data[4088]=0;
        data[4087]=0;
        data[4086]=0;
        data[4085]=0;
        data[4084]=0;
        data[4083]=0;
        data[4082]=0;
        data[4081]=0;
        data[4080]=0;
        data[4079]=0;
        data[4078]=0;
        data[4077]=0;
        data[4076]=0;
        data[4075]=0;
        data[4074]=0;
        data[4073]=0;
        data[4072]=0;
        data[4071]=0;
        data[4070]=3;
        data[4069]=5;
        data[4068]=8;
        data[4067]=10;
        data[4066]=13;
        data[4065]=15;
        data[4064]=18;
        data[4063]=20;
        data[4062]=23;
        data[4061]=25;
        data[4060]=28;
        data[4059]=31;
        data[4058]=33;
        data[4057]=36;
        data[4056]=38;
        data[4055]=41;
        data[4054]=43;
        data[4053]=46;
        data[4052]=48;
        data[4051]=51;
        data[4050]=54;
        data[4049]=56;
        data[4048]=59;
        data[4047]=61;
        data[4046]=64;
        data[4045]=66;
        data[4044]=69;
        data[4043]=71;
        data[4042]=74;
        data[4041]=77;
        data[4040]=79;
        data[4039]=82;
        data[4038]=84;
        data[4037]=87;
        data[4036]=89;
        data[4035]=92;
        data[4034]=94;
        data[4033]=97;
        data[4032]=99;
        data[4031]=102;
        data[4030]=105;
        data[4029]=107;
        data[4028]=110;
        data[4027]=112;
        data[4026]=115;
        data[4025]=117;
        data[4024]=120;
        data[4023]=122;
        data[4022]=125;
        data[4021]=127;
        data[4020]=130;
        data[4019]=133;
        data[4018]=135;
        data[4017]=138;
        data[4016]=140;
        data[4015]=143;
        data[4014]=145;
        data[4013]=148;
        data[4012]=150;
        data[4011]=153;
        data[4010]=156;
        data[4009]=158;
        data[4008]=161;
        data[4007]=163;
        data[4006]=166;
        data[4005]=168;
        data[4004]=171;
        data[4003]=173;
        data[4002]=176;
        data[4001]=179;
        data[4000]=181;
        data[3999]=184;
        data[3998]=186;
        data[3997]=189;
        data[3996]=191;
        data[3995]=194;
        data[3994]=196;
        data[3993]=199;
        data[3992]=201;
        data[3991]=204;
        data[3990]=207;
        data[3989]=209;
        data[3988]=212;
        data[3987]=214;
        data[3986]=217;
        data[3985]=219;
        data[3984]=222;
        data[3983]=224;
        data[3982]=227;
        data[3981]=229;
        data[3980]=232;
        data[3979]=235;
        data[3978]=237;
        data[3977]=240;
        data[3976]=242;
        data[3975]=245;
        data[3974]=247;
        data[3973]=250;
        data[3972]=252;
        data[3971]=255;
        data[3970]=254;
        data[3969]=254;
        data[3968]=254;
        data[3967]=254;
        data[3966]=253;
        data[3965]=253;
        data[3964]=253;
        data[3963]=252;
        data[3962]=252;
        data[3961]=252;
        data[3960]=252;
        data[3959]=251;
        data[3958]=251;
        data[3957]=251;
        data[3956]=250;
        data[3955]=250;
        data[3954]=250;
        data[3953]=250;
        data[3952]=249;
        data[3951]=249;
        data[3950]=249;
        data[3949]=248;
        data[3948]=248;
        data[3947]=248;
        data[3946]=248;
        data[3945]=247;
        data[3944]=247;
        data[3943]=247;
        data[3942]=247;
        data[3941]=246;
        data[3940]=246;
        data[3939]=246;
        data[3938]=245;
        data[3937]=245;
        data[3936]=245;
        data[3935]=245;
        data[3934]=244;
        data[3933]=244;
        data[3932]=244;
        data[3931]=243;
        data[3930]=243;
        data[3929]=243;
        data[3928]=243;
        data[3927]=242;
        data[3926]=242;
        data[3925]=242;
        data[3924]=241;
        data[3923]=241;
        data[3922]=241;
        data[3921]=241;
        data[3920]=240;
        data[3919]=240;
        data[3918]=240;
        data[3917]=239;
        data[3916]=239;
        data[3915]=239;
        data[3914]=239;
        data[3913]=238;
        data[3912]=238;
        data[3911]=238;
        data[3910]=237;
        data[3909]=237;
        data[3908]=237;
        data[3907]=237;
        data[3906]=236;
        data[3905]=236;
        data[3904]=236;
        data[3903]=235;
        data[3902]=235;
        data[3901]=235;
        data[3900]=235;
        data[3899]=234;
        data[3898]=234;
        data[3897]=234;
        data[3896]=233;
        data[3895]=233;
        data[3894]=233;
        data[3893]=233;
        data[3892]=232;
        data[3891]=232;
        data[3890]=232;
        data[3889]=231;
        data[3888]=231;
        data[3887]=231;
        data[3886]=231;
        data[3885]=230;
        data[3884]=230;
        data[3883]=230;
        data[3882]=229;
        data[3881]=229;
        data[3880]=229;
        data[3879]=229;
        data[3878]=228;
        data[3877]=228;
        data[3876]=228;
        data[3875]=228;
        data[3874]=227;
        data[3873]=227;
        data[3872]=227;
        data[3871]=226;
        data[3870]=226;
        data[3869]=226;
        data[3868]=226;
        data[3867]=225;
        data[3866]=225;
        data[3865]=225;
        data[3864]=224;
        data[3863]=224;
        data[3862]=224;
        data[3861]=224;
        data[3860]=223;
        data[3859]=223;
        data[3858]=223;
        data[3857]=222;
        data[3856]=222;
        data[3855]=222;
        data[3854]=222;
        data[3853]=221;
        data[3852]=221;
        data[3851]=221;
        data[3850]=220;
        data[3849]=220;
        data[3848]=220;
        data[3847]=220;
        data[3846]=219;
        data[3845]=219;
        data[3844]=219;
        data[3843]=218;
        data[3842]=218;
        data[3841]=218;
        data[3840]=218;
        data[3839]=217;
        data[3838]=217;
        data[3837]=217;
        data[3836]=216;
        data[3835]=216;
        data[3834]=216;
        data[3833]=216;
        data[3832]=215;
        data[3831]=215;
        data[3830]=215;
        data[3829]=214;
        data[3828]=214;
        data[3827]=214;
        data[3826]=214;
        data[3825]=213;
        data[3824]=213;
        data[3823]=213;
        data[3822]=213;
        data[3821]=212;
        data[3820]=212;
        data[3819]=212;
        data[3818]=211;
        data[3817]=211;
        data[3816]=211;
        data[3815]=211;
        data[3814]=210;
        data[3813]=210;
        data[3812]=210;
        data[3811]=209;
        data[3810]=209;
        data[3809]=209;
        data[3808]=209;
        data[3807]=208;
        data[3806]=208;
        data[3805]=208;
        data[3804]=207;
        data[3803]=207;
        data[3802]=207;
        data[3801]=207;
        data[3800]=206;
        data[3799]=206;
        data[3798]=206;
        data[3797]=205;
        data[3796]=205;
        data[3795]=205;
        data[3794]=205;
        data[3793]=204;
        data[3792]=204;
        data[3791]=204;
        data[3790]=203;
        data[3789]=203;
        data[3788]=203;
        data[3787]=203;
        data[3786]=202;
        data[3785]=202;
        data[3784]=202;
        data[3783]=201;
        data[3782]=201;
        data[3781]=201;
        data[3780]=201;
        data[3779]=200;
        data[3778]=200;
        data[3777]=200;
        data[3776]=199;
        data[3775]=199;
        data[3774]=199;
        data[3773]=199;
        data[3772]=198;
        data[3771]=198;
        data[3770]=198;
        data[3769]=197;
        data[3768]=197;
        data[3767]=197;
        data[3766]=197;
        data[3765]=196;
        data[3764]=196;
        data[3763]=196;
        data[3762]=195;
        data[3761]=195;
        data[3760]=195;
        data[3759]=195;
        data[3758]=194;
        data[3757]=194;
        data[3756]=194;
        data[3755]=194;
        data[3754]=193;
        data[3753]=193;
        data[3752]=193;
        data[3751]=192;
        data[3750]=192;
        data[3749]=192;
        data[3748]=192;
        data[3747]=191;
        data[3746]=191;
        data[3745]=191;
        data[3744]=190;
        data[3743]=190;
        data[3742]=190;
        data[3741]=190;
        data[3740]=189;
        data[3739]=189;
        data[3738]=189;
        data[3737]=188;
        data[3736]=188;
        data[3735]=188;
        data[3734]=188;
        data[3733]=187;
        data[3732]=187;
        data[3731]=187;
        data[3730]=186;
        data[3729]=186;
        data[3728]=186;
        data[3727]=186;
        data[3726]=185;
        data[3725]=185;
        data[3724]=185;
        data[3723]=184;
        data[3722]=184;
        data[3721]=184;
        data[3720]=184;
        data[3719]=183;
        data[3718]=183;
        data[3717]=183;
        data[3716]=182;
        data[3715]=182;
        data[3714]=182;
        data[3713]=182;
        data[3712]=181;
        data[3711]=181;
        data[3710]=181;
        data[3709]=180;
        data[3708]=180;
        data[3707]=180;
        data[3706]=180;
        data[3705]=179;
        data[3704]=179;
        data[3703]=179;
        data[3702]=178;
        data[3701]=178;
        data[3700]=178;
        data[3699]=178;
        data[3698]=177;
        data[3697]=177;
        data[3696]=177;
        data[3695]=177;
        data[3694]=176;
        data[3693]=176;
        data[3692]=176;
        data[3691]=175;
        data[3690]=175;
        data[3689]=175;
        data[3688]=175;
        data[3687]=174;
        data[3686]=174;
        data[3685]=174;
        data[3684]=173;
        data[3683]=173;
        data[3682]=173;
        data[3681]=173;
        data[3680]=172;
        data[3679]=172;
        data[3678]=172;
        data[3677]=171;
        data[3676]=171;
        data[3675]=171;
        data[3674]=171;
        data[3673]=170;
        data[3672]=170;
        data[3671]=170;
        data[3670]=169;
        data[3669]=169;
        data[3668]=169;
        data[3667]=169;
        data[3666]=168;
        data[3665]=168;
        data[3664]=168;
        data[3663]=167;
        data[3662]=167;
        data[3661]=167;
        data[3660]=167;
        data[3659]=166;
        data[3658]=166;
        data[3657]=166;
        data[3656]=165;
        data[3655]=165;
        data[3654]=165;
        data[3653]=165;
        data[3652]=164;
        data[3651]=164;
        data[3650]=164;
        data[3649]=163;
        data[3648]=163;
        data[3647]=163;
        data[3646]=163;
        data[3645]=162;
        data[3644]=162;
        data[3643]=162;
        data[3642]=162;
        data[3641]=161;
        data[3640]=161;
        data[3639]=161;
        data[3638]=160;
        data[3637]=160;
        data[3636]=160;
        data[3635]=160;
        data[3634]=159;
        data[3633]=159;
        data[3632]=159;
        data[3631]=158;
        data[3630]=158;
        data[3629]=158;
        data[3628]=158;
        data[3627]=157;
        data[3626]=157;
        data[3625]=157;
        data[3624]=156;
        data[3623]=156;
        data[3622]=156;
        data[3621]=156;
        data[3620]=155;
        data[3619]=155;
        data[3618]=155;
        data[3617]=154;
        data[3616]=154;
        data[3615]=154;
        data[3614]=154;
        data[3613]=153;
        data[3612]=153;
        data[3611]=153;
        data[3610]=152;
        data[3609]=152;
        data[3608]=152;
        data[3607]=152;
        data[3606]=151;
        data[3605]=151;
        data[3604]=151;
        data[3603]=150;
        data[3602]=150;
        data[3601]=150;
        data[3600]=150;
        data[3599]=149;
        data[3598]=149;
        data[3597]=149;
        data[3596]=148;
        data[3595]=148;
        data[3594]=148;
        data[3593]=148;
        data[3592]=147;
        data[3591]=147;
        data[3590]=147;
        data[3589]=146;
        data[3588]=146;
        data[3587]=146;
        data[3586]=146;
        data[3585]=145;
        data[3584]=145;
        data[3583]=145;
        data[3582]=144;
        data[3581]=144;
        data[3580]=144;
        data[3579]=144;
        data[3578]=143;
        data[3577]=143;
        data[3576]=143;
        data[3575]=143;
        data[3574]=142;
        data[3573]=142;
        data[3572]=142;
        data[3571]=141;
        data[3570]=141;
        data[3569]=141;
        data[3568]=141;
        data[3567]=140;
        data[3566]=140;
        data[3565]=140;
        data[3564]=139;
        data[3563]=139;
        data[3562]=139;
        data[3561]=139;
        data[3560]=138;
        data[3559]=138;
        data[3558]=138;
        data[3557]=137;
        data[3556]=137;
        data[3555]=137;
        data[3554]=137;
        data[3553]=136;
        data[3552]=136;
        data[3551]=136;
        data[3550]=135;
        data[3549]=135;
        data[3548]=135;
        data[3547]=135;
        data[3546]=134;
        data[3545]=134;
        data[3544]=134;
        data[3543]=133;
        data[3542]=133;
        data[3541]=133;
        data[3540]=133;
        data[3539]=132;
        data[3538]=132;
        data[3537]=132;
        data[3536]=131;
        data[3535]=131;
        data[3534]=131;
        data[3533]=131;
        data[3532]=130;
        data[3531]=130;
        data[3530]=130;
        data[3529]=129;
        data[3528]=129;
        data[3527]=129;
        data[3526]=129;
        data[3525]=128;
        data[3524]=128;
        data[3523]=128;
        data[3522]=128;
        data[3521]=127;
        data[3520]=127;
        data[3519]=127;
        data[3518]=126;
        data[3517]=126;
        data[3516]=126;
        data[3515]=126;
        data[3514]=125;
        data[3513]=125;
        data[3512]=125;
        data[3511]=124;
        data[3510]=124;
        data[3509]=124;
        data[3508]=124;
        data[3507]=123;
        data[3506]=123;
        data[3505]=123;
        data[3504]=122;
        data[3503]=122;
        data[3502]=122;
        data[3501]=122;
        data[3500]=121;
        data[3499]=121;
        data[3498]=121;
        data[3497]=120;
        data[3496]=120;
        data[3495]=120;
        data[3494]=120;
        data[3493]=119;
        data[3492]=119;
        data[3491]=119;
        data[3490]=118;
        data[3489]=118;
        data[3488]=118;
        data[3487]=118;
        data[3486]=117;
        data[3485]=117;
        data[3484]=117;
        data[3483]=116;
        data[3482]=116;
        data[3481]=116;
        data[3480]=116;
        data[3479]=115;
        data[3478]=115;
        data[3477]=115;
        data[3476]=114;
        data[3475]=114;
        data[3474]=114;
        data[3473]=114;
        data[3472]=113;
        data[3471]=113;
        data[3470]=113;
        data[3469]=112;
        data[3468]=112;
        data[3467]=112;
        data[3466]=112;
        data[3465]=111;
        data[3464]=111;
        data[3463]=111;
        data[3462]=110;
        data[3461]=110;
        data[3460]=110;
        data[3459]=110;
        data[3458]=109;
        data[3457]=109;
        data[3456]=109;
        data[3455]=109;
        data[3454]=108;
        data[3453]=108;
        data[3452]=108;
        data[3451]=107;
        data[3450]=107;
        data[3449]=107;
        data[3448]=107;
        data[3447]=106;
        data[3446]=106;
        data[3445]=106;
        data[3444]=105;
        data[3443]=105;
        data[3442]=105;
        data[3441]=105;
        data[3440]=104;
        data[3439]=104;
        data[3438]=104;
        data[3437]=103;
        data[3436]=103;
        data[3435]=103;
        data[3434]=103;
        data[3433]=102;
        data[3432]=102;
        data[3431]=102;
        data[3430]=101;
        data[3429]=101;
        data[3428]=101;
        data[3427]=101;
        data[3426]=100;
        data[3425]=100;
        data[3424]=100;
        data[3423]=99;
        data[3422]=99;
        data[3421]=99;
        data[3420]=99;
        data[3419]=98;
        data[3418]=98;
        data[3417]=98;
        data[3416]=97;
        data[3415]=97;
        data[3414]=97;
        data[3413]=97;
        data[3412]=96;
        data[3411]=96;
        data[3410]=96;
        data[3409]=95;
        data[3408]=95;
        data[3407]=95;
        data[3406]=95;
        data[3405]=94;
        data[3404]=94;
        data[3403]=94;
        data[3402]=94;
        data[3401]=93;
        data[3400]=93;
        data[3399]=93;
        data[3398]=92;
        data[3397]=92;
        data[3396]=92;
        data[3395]=92;
        data[3394]=91;
        data[3393]=91;
        data[3392]=91;
        data[3391]=90;
        data[3390]=90;
        data[3389]=90;
        data[3388]=90;
        data[3387]=89;
        data[3386]=89;
        data[3385]=89;
        data[3384]=88;
        data[3383]=88;
        data[3382]=88;
        data[3381]=88;
        data[3380]=87;
        data[3379]=87;
        data[3378]=87;
        data[3377]=86;
        data[3376]=86;
        data[3375]=86;
        data[3374]=86;
        data[3373]=85;
        data[3372]=85;
        data[3371]=85;
        data[3370]=84;
        data[3369]=84;
        data[3368]=84;
        data[3367]=84;
        data[3366]=83;
        data[3365]=83;
        data[3364]=83;
        data[3363]=82;
        data[3362]=82;
        data[3361]=82;
        data[3360]=82;
        data[3359]=81;
        data[3358]=81;
        data[3357]=81;
        data[3356]=80;
        data[3355]=80;
        data[3354]=80;
        data[3353]=80;
        data[3352]=79;
        data[3351]=79;
        data[3350]=79;
        data[3349]=78;
        data[3348]=78;
        data[3347]=78;
        data[3346]=78;
        data[3345]=77;
        data[3344]=77;
        data[3343]=77;
        data[3342]=77;
        data[3341]=76;
        data[3340]=76;
        data[3339]=76;
        data[3338]=75;
        data[3337]=75;
        data[3336]=75;
        data[3335]=75;
        data[3334]=74;
        data[3333]=74;
        data[3332]=74;
        data[3331]=73;
        data[3330]=73;
        data[3329]=73;
        data[3328]=73;
        data[3327]=72;
        data[3326]=72;
        data[3325]=72;
        data[3324]=71;
        data[3323]=71;
        data[3322]=71;
        data[3321]=71;
        data[3320]=70;
        data[3319]=70;
        data[3318]=70;
        data[3317]=69;
        data[3316]=69;
        data[3315]=69;
        data[3314]=69;
        data[3313]=68;
        data[3312]=68;
        data[3311]=68;
        data[3310]=67;
        data[3309]=67;
        data[3308]=67;
        data[3307]=67;
        data[3306]=66;
        data[3305]=66;
        data[3304]=66;
        data[3303]=65;
        data[3302]=65;
        data[3301]=65;
        data[3300]=65;
        data[3299]=64;
        data[3298]=64;
        data[3297]=64;
        data[3296]=63;
        data[3295]=63;
        data[3294]=63;
        data[3293]=63;
        data[3292]=62;
        data[3291]=62;
        data[3290]=62;
        data[3289]=61;
        data[3288]=61;
        data[3287]=61;
        data[3286]=61;
        data[3285]=60;
        data[3284]=60;
        data[3283]=60;
        data[3282]=59;
        data[3281]=59;
        data[3280]=59;
        data[3279]=59;
        data[3278]=58;
        data[3277]=58;
        data[3276]=58;
        data[3275]=58;
        data[3274]=57;
        data[3273]=57;
        data[3272]=57;
        data[3271]=56;
        data[3270]=56;
        data[3269]=56;
        data[3268]=56;
        data[3267]=55;
        data[3266]=55;
        data[3265]=55;
        data[3264]=54;
        data[3263]=54;
        data[3262]=54;
        data[3261]=54;
        data[3260]=53;
        data[3259]=53;
        data[3258]=53;
        data[3257]=52;
        data[3256]=52;
        data[3255]=52;
        data[3254]=52;
        data[3253]=51;
        data[3252]=51;
        data[3251]=51;
        data[3250]=50;
        data[3249]=50;
        data[3248]=50;
        data[3247]=50;
        data[3246]=49;
        data[3245]=49;
        data[3244]=49;
        data[3243]=48;
        data[3242]=48;
        data[3241]=48;
        data[3240]=48;
        data[3239]=47;
        data[3238]=47;
        data[3237]=47;
        data[3236]=46;
        data[3235]=46;
        data[3234]=46;
        data[3233]=46;
        data[3232]=45;
        data[3231]=45;
        data[3230]=45;
        data[3229]=44;
        data[3228]=44;
        data[3227]=44;
        data[3226]=44;
        data[3225]=43;
        data[3224]=43;
        data[3223]=43;
        data[3222]=43;
        data[3221]=42;
        data[3220]=42;
        data[3219]=42;
        data[3218]=41;
        data[3217]=41;
        data[3216]=41;
        data[3215]=41;
        data[3214]=40;
        data[3213]=40;
        data[3212]=40;
        data[3211]=39;
        data[3210]=39;
        data[3209]=39;
        data[3208]=39;
        data[3207]=38;
        data[3206]=38;
        data[3205]=38;
        data[3204]=37;
        data[3203]=37;
        data[3202]=37;
        data[3201]=37;
        data[3200]=36;
        data[3199]=36;
        data[3198]=36;
        data[3197]=35;
        data[3196]=35;
        data[3195]=35;
        data[3194]=35;
        data[3193]=34;
        data[3192]=34;
        data[3191]=34;
        data[3190]=33;
        data[3189]=33;
        data[3188]=33;
        data[3187]=33;
        data[3186]=32;
        data[3185]=32;
        data[3184]=32;
        data[3183]=31;
        data[3182]=31;
        data[3181]=31;
        data[3180]=31;
        data[3179]=30;
        data[3178]=30;
        data[3177]=30;
        data[3176]=29;
        data[3175]=29;
        data[3174]=29;
        data[3173]=29;
        data[3172]=28;
        data[3171]=28;
        data[3170]=28;
        data[3169]=27;
        data[3168]=27;
        data[3167]=27;
        data[3166]=27;
        data[3165]=26;
        data[3164]=26;
        data[3163]=26;
        data[3162]=25;
        data[3161]=25;
        data[3160]=25;
        data[3159]=25;
        data[3158]=24;
        data[3157]=24;
        data[3156]=24;
        data[3155]=24;
        data[3154]=23;
        data[3153]=23;
        data[3152]=23;
        data[3151]=22;
        data[3150]=22;
        data[3149]=22;
        data[3148]=22;
        data[3147]=21;
        data[3146]=21;
        data[3145]=21;
        data[3144]=20;
        data[3143]=20;
        data[3142]=20;
        data[3141]=20;
        data[3140]=19;
        data[3139]=19;
        data[3138]=19;
        data[3137]=18;
        data[3136]=18;
        data[3135]=18;
        data[3134]=18;
        data[3133]=17;
        data[3132]=17;
        data[3131]=17;
        data[3130]=16;
        data[3129]=16;
        data[3128]=16;
        data[3127]=16;
        data[3126]=15;
        data[3125]=15;
        data[3124]=15;
        data[3123]=14;
        data[3122]=14;
        data[3121]=14;
        data[3120]=14;
        data[3119]=13;
        data[3118]=13;
        data[3117]=13;
        data[3116]=12;
        data[3115]=12;
        data[3114]=12;
        data[3113]=12;
        data[3112]=11;
        data[3111]=11;
        data[3110]=11;
        data[3109]=10;
        data[3108]=10;
        data[3107]=10;
        data[3106]=10;
        data[3105]=9;
        data[3104]=9;
        data[3103]=9;
        data[3102]=9;
        data[3101]=8;
        data[3100]=8;
        data[3099]=8;
        data[3098]=7;
        data[3097]=7;
        data[3096]=7;
        data[3095]=7;
        data[3094]=6;
        data[3093]=6;
        data[3092]=6;
        data[3091]=5;
        data[3090]=5;
        data[3089]=5;
        data[3088]=5;
        data[3087]=4;
        data[3086]=4;
        data[3085]=4;
        data[3084]=3;
        data[3083]=3;
        data[3082]=3;
        data[3081]=3;
        data[3080]=2;
        data[3079]=2;
        data[3078]=2;
        data[3077]=1;
        data[3076]=1;
        data[3075]=1;
        data[3074]=1;
        data[3073]=0;
        data[3072]=0;
        data[3071]=0;
        data[3070]=0;
        data[3069]=0;
        data[3068]=0;
        data[3067]=0;
        data[3066]=0;
        data[3065]=0;
        data[3064]=0;
        data[3063]=0;
        data[3062]=0;
        data[3061]=0;
        data[3060]=0;
        data[3059]=0;
        data[3058]=0;
        data[3057]=0;
        data[3056]=0;
        data[3055]=0;
        data[3054]=0;
        data[3053]=0;
        data[3052]=0;
        data[3051]=0;
        data[3050]=0;
        data[3049]=0;
        data[3048]=0;
        data[3047]=0;
        data[3046]=1;
        data[3045]=1;
        data[3044]=2;
        data[3043]=2;
        data[3042]=3;
        data[3041]=3;
        data[3040]=4;
        data[3039]=4;
        data[3038]=5;
        data[3037]=5;
        data[3036]=6;
        data[3035]=6;
        data[3034]=7;
        data[3033]=7;
        data[3032]=8;
        data[3031]=8;
        data[3030]=9;
        data[3029]=9;
        data[3028]=10;
        data[3027]=10;
        data[3026]=11;
        data[3025]=11;
        data[3024]=12;
        data[3023]=12;
        data[3022]=13;
        data[3021]=13;
        data[3020]=14;
        data[3019]=14;
        data[3018]=15;
        data[3017]=15;
        data[3016]=16;
        data[3015]=16;
        data[3014]=17;
        data[3013]=17;
        data[3012]=18;
        data[3011]=18;
        data[3010]=19;
        data[3009]=19;
        data[3008]=20;
        data[3007]=20;
        data[3006]=21;
        data[3005]=21;
        data[3004]=22;
        data[3003]=22;
        data[3002]=23;
        data[3001]=23;
        data[3000]=24;
        data[2999]=24;
        data[2998]=25;
        data[2997]=25;
        data[2996]=26;
        data[2995]=27;
        data[2994]=27;
        data[2993]=28;
        data[2992]=28;
        data[2991]=29;
        data[2990]=29;
        data[2989]=30;
        data[2988]=30;
        data[2987]=31;
        data[2986]=31;
        data[2985]=32;
        data[2984]=32;
        data[2983]=33;
        data[2982]=33;
        data[2981]=34;
        data[2980]=34;
        data[2979]=35;
        data[2978]=35;
        data[2977]=36;
        data[2976]=36;
        data[2975]=37;
        data[2974]=37;
        data[2973]=38;
        data[2972]=38;
        data[2971]=39;
        data[2970]=39;
        data[2969]=40;
        data[2968]=40;
        data[2967]=41;
        data[2966]=41;
        data[2965]=42;
        data[2964]=42;
        data[2963]=43;
        data[2962]=43;
        data[2961]=44;
        data[2960]=44;
        data[2959]=45;
        data[2958]=45;
        data[2957]=46;
        data[2956]=46;
        data[2955]=47;
        data[2954]=47;
        data[2953]=48;
        data[2952]=48;
        data[2951]=49;
        data[2950]=49;
        data[2949]=50;
        data[2948]=50;
        data[2947]=51;
        data[2946]=52;
        data[2945]=52;
        data[2944]=53;
        data[2943]=53;
        data[2942]=54;
        data[2941]=54;
        data[2940]=55;
        data[2939]=55;
        data[2938]=56;
        data[2937]=56;
        data[2936]=57;
        data[2935]=57;
        data[2934]=58;
        data[2933]=58;
        data[2932]=59;
        data[2931]=59;
        data[2930]=60;
        data[2929]=60;
        data[2928]=61;
        data[2927]=61;
        data[2926]=62;
        data[2925]=62;
        data[2924]=63;
        data[2923]=63;
        data[2922]=64;
        data[2921]=64;
        data[2920]=65;
        data[2919]=65;
        data[2918]=66;
        data[2917]=66;
        data[2916]=67;
        data[2915]=67;
        data[2914]=68;
        data[2913]=68;
        data[2912]=69;
        data[2911]=69;
        data[2910]=70;
        data[2909]=70;
        data[2908]=71;
        data[2907]=71;
        data[2906]=72;
        data[2905]=72;
        data[2904]=73;
        data[2903]=73;
        data[2902]=74;
        data[2901]=74;
        data[2900]=75;
        data[2899]=75;
        data[2898]=76;
        data[2897]=77;
        data[2896]=77;
        data[2895]=78;
        data[2894]=78;
        data[2893]=79;
        data[2892]=79;
        data[2891]=80;
        data[2890]=80;
        data[2889]=81;
        data[2888]=81;
        data[2887]=82;
        data[2886]=82;
        data[2885]=83;
        data[2884]=83;
        data[2883]=84;
        data[2882]=84;
        data[2881]=85;
        data[2880]=85;
        data[2879]=86;
        data[2878]=86;
        data[2877]=87;
        data[2876]=87;
        data[2875]=88;
        data[2874]=88;
        data[2873]=89;
        data[2872]=89;
        data[2871]=90;
        data[2870]=90;
        data[2869]=91;
        data[2868]=91;
        data[2867]=92;
        data[2866]=92;
        data[2865]=93;
        data[2864]=93;
        data[2863]=94;
        data[2862]=94;
        data[2861]=95;
        data[2860]=95;
        data[2859]=96;
        data[2858]=96;
        data[2857]=97;
        data[2856]=97;
        data[2855]=98;
        data[2854]=98;
        data[2853]=99;
        data[2852]=99;
        data[2851]=100;
        data[2850]=100;
        data[2849]=101;
        data[2848]=101;
        data[2847]=102;
        data[2846]=103;
        data[2845]=103;
        data[2844]=104;
        data[2843]=104;
        data[2842]=105;
        data[2841]=105;
        data[2840]=106;
        data[2839]=106;
        data[2838]=107;
        data[2837]=107;
        data[2836]=108;
        data[2835]=108;
        data[2834]=109;
        data[2833]=109;
        data[2832]=110;
        data[2831]=110;
        data[2830]=111;
        data[2829]=111;
        data[2828]=112;
        data[2827]=112;
        data[2826]=113;
        data[2825]=113;
        data[2824]=114;
        data[2823]=114;
        data[2822]=115;
        data[2821]=115;
        data[2820]=116;
        data[2819]=116;
        data[2818]=117;
        data[2817]=117;
        data[2816]=118;
        data[2815]=118;
        data[2814]=119;
        data[2813]=119;
        data[2812]=120;
        data[2811]=120;
        data[2810]=121;
        data[2809]=121;
        data[2808]=122;
        data[2807]=122;
        data[2806]=123;
        data[2805]=123;
        data[2804]=124;
        data[2803]=124;
        data[2802]=125;
        data[2801]=125;
        data[2800]=126;
        data[2799]=126;
        data[2798]=127;
        data[2797]=128;
        data[2796]=128;
        data[2795]=129;
        data[2794]=129;
        data[2793]=130;
        data[2792]=130;
        data[2791]=131;
        data[2790]=131;
        data[2789]=132;
        data[2788]=132;
        data[2787]=133;
        data[2786]=133;
        data[2785]=134;
        data[2784]=134;
        data[2783]=135;
        data[2782]=135;
        data[2781]=136;
        data[2780]=136;
        data[2779]=137;
        data[2778]=137;
        data[2777]=138;
        data[2776]=138;
        data[2775]=139;
        data[2774]=139;
        data[2773]=140;
        data[2772]=140;
        data[2771]=141;
        data[2770]=141;
        data[2769]=142;
        data[2768]=142;
        data[2767]=143;
        data[2766]=143;
        data[2765]=144;
        data[2764]=144;
        data[2763]=145;
        data[2762]=145;
        data[2761]=146;
        data[2760]=146;
        data[2759]=147;
        data[2758]=147;
        data[2757]=148;
        data[2756]=148;
        data[2755]=149;
        data[2754]=149;
        data[2753]=150;
        data[2752]=150;
        data[2751]=151;
        data[2750]=151;
        data[2749]=152;
        data[2748]=152;
        data[2747]=153;
        data[2746]=154;
        data[2745]=154;
        data[2744]=155;
        data[2743]=155;
        data[2742]=156;
        data[2741]=156;
        data[2740]=157;
        data[2739]=157;
        data[2738]=158;
        data[2737]=158;
        data[2736]=159;
        data[2735]=159;
        data[2734]=160;
        data[2733]=160;
        data[2732]=161;
        data[2731]=161;
        data[2730]=162;
        data[2729]=162;
        data[2728]=163;
        data[2727]=163;
        data[2726]=164;
        data[2725]=164;
        data[2724]=165;
        data[2723]=165;
        data[2722]=166;
        data[2721]=166;
        data[2720]=167;
        data[2719]=167;
        data[2718]=168;
        data[2717]=168;
        data[2716]=169;
        data[2715]=169;
        data[2714]=170;
        data[2713]=170;
        data[2712]=171;
        data[2711]=171;
        data[2710]=172;
        data[2709]=172;
        data[2708]=173;
        data[2707]=173;
        data[2706]=174;
        data[2705]=174;
        data[2704]=175;
        data[2703]=175;
        data[2702]=176;
        data[2701]=176;
        data[2700]=177;
        data[2699]=177;
        data[2698]=178;
        data[2697]=179;
        data[2696]=179;
        data[2695]=180;
        data[2694]=180;
        data[2693]=181;
        data[2692]=181;
        data[2691]=182;
        data[2690]=182;
        data[2689]=183;
        data[2688]=183;
        data[2687]=184;
        data[2686]=184;
        data[2685]=185;
        data[2684]=185;
        data[2683]=186;
        data[2682]=186;
        data[2681]=187;
        data[2680]=187;
        data[2679]=188;
        data[2678]=188;
        data[2677]=189;
        data[2676]=189;
        data[2675]=190;
        data[2674]=190;
        data[2673]=191;
        data[2672]=191;
        data[2671]=192;
        data[2670]=192;
        data[2669]=193;
        data[2668]=193;
        data[2667]=194;
        data[2666]=194;
        data[2665]=195;
        data[2664]=195;
        data[2663]=196;
        data[2662]=196;
        data[2661]=197;
        data[2660]=197;
        data[2659]=198;
        data[2658]=198;
        data[2657]=199;
        data[2656]=199;
        data[2655]=200;
        data[2654]=200;
        data[2653]=201;
        data[2652]=201;
        data[2651]=202;
        data[2650]=202;
        data[2649]=203;
        data[2648]=203;
        data[2647]=204;
        data[2646]=205;
        data[2645]=205;
        data[2644]=206;
        data[2643]=206;
        data[2642]=207;
        data[2641]=207;
        data[2640]=208;
        data[2639]=208;
        data[2638]=209;
        data[2637]=209;
        data[2636]=210;
        data[2635]=210;
        data[2634]=211;
        data[2633]=211;
        data[2632]=212;
        data[2631]=212;
        data[2630]=213;
        data[2629]=213;
        data[2628]=214;
        data[2627]=214;
        data[2626]=215;
        data[2625]=215;
        data[2624]=216;
        data[2623]=216;
        data[2622]=217;
        data[2621]=217;
        data[2620]=218;
        data[2619]=218;
        data[2618]=219;
        data[2617]=219;
        data[2616]=220;
        data[2615]=220;
        data[2614]=221;
        data[2613]=221;
        data[2612]=222;
        data[2611]=222;
        data[2610]=223;
        data[2609]=223;
        data[2608]=224;
        data[2607]=224;
        data[2606]=225;
        data[2605]=225;
        data[2604]=226;
        data[2603]=226;
        data[2602]=227;
        data[2601]=227;
        data[2600]=228;
        data[2599]=228;
        data[2598]=229;
        data[2597]=230;
        data[2596]=230;
        data[2595]=231;
        data[2594]=231;
        data[2593]=232;
        data[2592]=232;
        data[2591]=233;
        data[2590]=233;
        data[2589]=234;
        data[2588]=234;
        data[2587]=235;
        data[2586]=235;
        data[2585]=236;
        data[2584]=236;
        data[2583]=237;
        data[2582]=237;
        data[2581]=238;
        data[2580]=238;
        data[2579]=239;
        data[2578]=239;
        data[2577]=240;
        data[2576]=240;
        data[2575]=241;
        data[2574]=241;
        data[2573]=242;
        data[2572]=242;
        data[2571]=243;
        data[2570]=243;
        data[2569]=244;
        data[2568]=244;
        data[2567]=245;
        data[2566]=245;
        data[2565]=246;
        data[2564]=246;
        data[2563]=247;
        data[2562]=247;
        data[2561]=248;
        data[2560]=248;
        data[2559]=249;
        data[2558]=249;
        data[2557]=250;
        data[2556]=250;
        data[2555]=251;
        data[2554]=251;
        data[2553]=252;
        data[2552]=252;
        data[2551]=253;
        data[2550]=253;
        data[2549]=254;
        data[2548]=254;
        data[2547]=254;
        data[2546]=254;
        data[2545]=253;
        data[2544]=253;
        data[2543]=252;
        data[2542]=252;
        data[2541]=251;
        data[2540]=251;
        data[2539]=250;
        data[2538]=250;
        data[2537]=249;
        data[2536]=249;
        data[2535]=248;
        data[2534]=248;
        data[2533]=247;
        data[2532]=247;
        data[2531]=246;
        data[2530]=246;
        data[2529]=245;
        data[2528]=245;
        data[2527]=244;
        data[2526]=244;
        data[2525]=243;
        data[2524]=243;
        data[2523]=242;
        data[2522]=242;
        data[2521]=241;
        data[2520]=241;
        data[2519]=240;
        data[2518]=240;
        data[2517]=239;
        data[2516]=239;
        data[2515]=238;
        data[2514]=238;
        data[2513]=237;
        data[2512]=237;
        data[2511]=236;
        data[2510]=236;
        data[2509]=235;
        data[2508]=235;
        data[2507]=234;
        data[2506]=234;
        data[2505]=233;
        data[2504]=233;
        data[2503]=232;
        data[2502]=232;
        data[2501]=231;
        data[2500]=231;
        data[2499]=230;
        data[2498]=230;
        data[2497]=229;
        data[2496]=228;
        data[2495]=228;
        data[2494]=227;
        data[2493]=227;
        data[2492]=226;
        data[2491]=226;
        data[2490]=225;
        data[2489]=225;
        data[2488]=224;
        data[2487]=224;
        data[2486]=223;
        data[2485]=223;
        data[2484]=222;
        data[2483]=222;
        data[2482]=221;
        data[2481]=221;
        data[2480]=220;
        data[2479]=220;
        data[2478]=219;
        data[2477]=219;
        data[2476]=218;
        data[2475]=218;
        data[2474]=217;
        data[2473]=217;
        data[2472]=216;
        data[2471]=216;
        data[2470]=215;
        data[2469]=215;
        data[2468]=214;
        data[2467]=214;
        data[2466]=213;
        data[2465]=213;
        data[2464]=212;
        data[2463]=212;
        data[2462]=211;
        data[2461]=211;
        data[2460]=210;
        data[2459]=210;
        data[2458]=209;
        data[2457]=209;
        data[2456]=208;
        data[2455]=208;
        data[2454]=207;
        data[2453]=207;
        data[2452]=206;
        data[2451]=206;
        data[2450]=205;
        data[2449]=205;
        data[2448]=204;
        data[2447]=203;
        data[2446]=203;
        data[2445]=202;
        data[2444]=202;
        data[2443]=201;
        data[2442]=201;
        data[2441]=200;
        data[2440]=200;
        data[2439]=199;
        data[2438]=199;
        data[2437]=198;
        data[2436]=198;
        data[2435]=197;
        data[2434]=197;
        data[2433]=196;
        data[2432]=196;
        data[2431]=195;
        data[2430]=195;
        data[2429]=194;
        data[2428]=194;
        data[2427]=193;
        data[2426]=193;
        data[2425]=192;
        data[2424]=192;
        data[2423]=191;
        data[2422]=191;
        data[2421]=190;
        data[2420]=190;
        data[2419]=189;
        data[2418]=189;
        data[2417]=188;
        data[2416]=188;
        data[2415]=187;
        data[2414]=187;
        data[2413]=186;
        data[2412]=186;
        data[2411]=185;
        data[2410]=185;
        data[2409]=184;
        data[2408]=184;
        data[2407]=183;
        data[2406]=183;
        data[2405]=182;
        data[2404]=182;
        data[2403]=181;
        data[2402]=181;
        data[2401]=180;
        data[2400]=180;
        data[2399]=179;
        data[2398]=179;
        data[2397]=178;
        data[2396]=177;
        data[2395]=177;
        data[2394]=176;
        data[2393]=176;
        data[2392]=175;
        data[2391]=175;
        data[2390]=174;
        data[2389]=174;
        data[2388]=173;
        data[2387]=173;
        data[2386]=172;
        data[2385]=172;
        data[2384]=171;
        data[2383]=171;
        data[2382]=170;
        data[2381]=170;
        data[2380]=169;
        data[2379]=169;
        data[2378]=168;
        data[2377]=168;
        data[2376]=167;
        data[2375]=167;
        data[2374]=166;
        data[2373]=166;
        data[2372]=165;
        data[2371]=165;
        data[2370]=164;
        data[2369]=164;
        data[2368]=163;
        data[2367]=163;
        data[2366]=162;
        data[2365]=162;
        data[2364]=161;
        data[2363]=161;
        data[2362]=160;
        data[2361]=160;
        data[2360]=159;
        data[2359]=159;
        data[2358]=158;
        data[2357]=158;
        data[2356]=157;
        data[2355]=157;
        data[2354]=156;
        data[2353]=156;
        data[2352]=155;
        data[2351]=155;
        data[2350]=154;
        data[2349]=154;
        data[2348]=153;
        data[2347]=152;
        data[2346]=152;
        data[2345]=151;
        data[2344]=151;
        data[2343]=150;
        data[2342]=150;
        data[2341]=149;
        data[2340]=149;
        data[2339]=148;
        data[2338]=148;
        data[2337]=147;
        data[2336]=147;
        data[2335]=146;
        data[2334]=146;
        data[2333]=145;
        data[2332]=145;
        data[2331]=144;
        data[2330]=144;
        data[2329]=143;
        data[2328]=143;
        data[2327]=142;
        data[2326]=142;
        data[2325]=141;
        data[2324]=141;
        data[2323]=140;
        data[2322]=140;
        data[2321]=139;
        data[2320]=139;
        data[2319]=138;
        data[2318]=138;
        data[2317]=137;
        data[2316]=137;
        data[2315]=136;
        data[2314]=136;
        data[2313]=135;
        data[2312]=135;
        data[2311]=134;
        data[2310]=134;
        data[2309]=133;
        data[2308]=133;
        data[2307]=132;
        data[2306]=132;
        data[2305]=131;
        data[2304]=131;
        data[2303]=130;
        data[2302]=130;
        data[2301]=129;
        data[2300]=129;
        data[2299]=128;
        data[2298]=128;
        data[2297]=127;
        data[2296]=126;
        data[2295]=126;
        data[2294]=125;
        data[2293]=125;
        data[2292]=124;
        data[2291]=124;
        data[2290]=123;
        data[2289]=123;
        data[2288]=122;
        data[2287]=122;
        data[2286]=121;
        data[2285]=121;
        data[2284]=120;
        data[2283]=120;
        data[2282]=119;
        data[2281]=119;
        data[2280]=118;
        data[2279]=118;
        data[2278]=117;
        data[2277]=117;
        data[2276]=116;
        data[2275]=116;
        data[2274]=115;
        data[2273]=115;
        data[2272]=114;
        data[2271]=114;
        data[2270]=113;
        data[2269]=113;
        data[2268]=112;
        data[2267]=112;
        data[2266]=111;
        data[2265]=111;
        data[2264]=110;
        data[2263]=110;
        data[2262]=109;
        data[2261]=109;
        data[2260]=108;
        data[2259]=108;
        data[2258]=107;
        data[2257]=107;
        data[2256]=106;
        data[2255]=106;
        data[2254]=105;
        data[2253]=105;
        data[2252]=104;
        data[2251]=104;
        data[2250]=103;
        data[2249]=103;
        data[2248]=102;
        data[2247]=101;
        data[2246]=101;
        data[2245]=100;
        data[2244]=100;
        data[2243]=99;
        data[2242]=99;
        data[2241]=98;
        data[2240]=98;
        data[2239]=97;
        data[2238]=97;
        data[2237]=96;
        data[2236]=96;
        data[2235]=95;
        data[2234]=95;
        data[2233]=94;
        data[2232]=94;
        data[2231]=93;
        data[2230]=93;
        data[2229]=92;
        data[2228]=92;
        data[2227]=91;
        data[2226]=91;
        data[2225]=90;
        data[2224]=90;
        data[2223]=89;
        data[2222]=89;
        data[2221]=88;
        data[2220]=88;
        data[2219]=87;
        data[2218]=87;
        data[2217]=86;
        data[2216]=86;
        data[2215]=85;
        data[2214]=85;
        data[2213]=84;
        data[2212]=84;
        data[2211]=83;
        data[2210]=83;
        data[2209]=82;
        data[2208]=82;
        data[2207]=81;
        data[2206]=81;
        data[2205]=80;
        data[2204]=80;
        data[2203]=79;
        data[2202]=79;
        data[2201]=78;
        data[2200]=78;
        data[2199]=77;
        data[2198]=77;
        data[2197]=76;
        data[2196]=75;
        data[2195]=75;
        data[2194]=74;
        data[2193]=74;
        data[2192]=73;
        data[2191]=73;
        data[2190]=72;
        data[2189]=72;
        data[2188]=71;
        data[2187]=71;
        data[2186]=70;
        data[2185]=70;
        data[2184]=69;
        data[2183]=69;
        data[2182]=68;
        data[2181]=68;
        data[2180]=67;
        data[2179]=67;
        data[2178]=66;
        data[2177]=66;
        data[2176]=65;
        data[2175]=65;
        data[2174]=64;
        data[2173]=64;
        data[2172]=63;
        data[2171]=63;
        data[2170]=62;
        data[2169]=62;
        data[2168]=61;
        data[2167]=61;
        data[2166]=60;
        data[2165]=60;
        data[2164]=59;
        data[2163]=59;
        data[2162]=58;
        data[2161]=58;
        data[2160]=57;
        data[2159]=57;
        data[2158]=56;
        data[2157]=56;
        data[2156]=55;
        data[2155]=55;
        data[2154]=54;
        data[2153]=54;
        data[2152]=53;
        data[2151]=53;
        data[2150]=52;
        data[2149]=52;
        data[2148]=51;
        data[2147]=50;
        data[2146]=50;
        data[2145]=49;
        data[2144]=49;
        data[2143]=48;
        data[2142]=48;
        data[2141]=47;
        data[2140]=47;
        data[2139]=46;
        data[2138]=46;
        data[2137]=45;
        data[2136]=45;
        data[2135]=44;
        data[2134]=44;
        data[2133]=43;
        data[2132]=43;
        data[2131]=42;
        data[2130]=42;
        data[2129]=41;
        data[2128]=41;
        data[2127]=40;
        data[2126]=40;
        data[2125]=39;
        data[2124]=39;
        data[2123]=38;
        data[2122]=38;
        data[2121]=37;
        data[2120]=37;
        data[2119]=36;
        data[2118]=36;
        data[2117]=35;
        data[2116]=35;
        data[2115]=34;
        data[2114]=34;
        data[2113]=33;
        data[2112]=33;
        data[2111]=32;
        data[2110]=32;
        data[2109]=31;
        data[2108]=31;
        data[2107]=30;
        data[2106]=30;
        data[2105]=29;
        data[2104]=29;
        data[2103]=28;
        data[2102]=28;
        data[2101]=27;
        data[2100]=27;
        data[2099]=26;
        data[2098]=25;
        data[2097]=25;
        data[2096]=24;
        data[2095]=24;
        data[2094]=23;
        data[2093]=23;
        data[2092]=22;
        data[2091]=22;
        data[2090]=21;
        data[2089]=21;
        data[2088]=20;
        data[2087]=20;
        data[2086]=19;
        data[2085]=19;
        data[2084]=18;
        data[2083]=18;
        data[2082]=17;
        data[2081]=17;
        data[2080]=16;
        data[2079]=16;
        data[2078]=15;
        data[2077]=15;
        data[2076]=14;
        data[2075]=14;
        data[2074]=13;
        data[2073]=13;
        data[2072]=12;
        data[2071]=12;
        data[2070]=11;
        data[2069]=11;
        data[2068]=10;
        data[2067]=10;
        data[2066]=9;
        data[2065]=9;
        data[2064]=8;
        data[2063]=8;
        data[2062]=7;
        data[2061]=7;
        data[2060]=6;
        data[2059]=6;
        data[2058]=5;
        data[2057]=5;
        data[2056]=4;
        data[2055]=4;
        data[2054]=3;
        data[2053]=3;
        data[2052]=2;
        data[2051]=2;
        data[2050]=1;
        data[2049]=1;
        data[2048]=0;
        data[2047]=0;
        data[2046]=0;
        data[2045]=0;
        data[2044]=0;
        data[2043]=0;
        data[2042]=0;
        data[2041]=0;
        data[2040]=0;
        data[2039]=0;
        data[2038]=0;
        data[2037]=0;
        data[2036]=0;
        data[2035]=0;
        data[2034]=0;
        data[2033]=0;
        data[2032]=0;
        data[2031]=0;
        data[2030]=0;
        data[2029]=0;
        data[2028]=0;
        data[2027]=0;
        data[2026]=0;
        data[2025]=0;
        data[2024]=0;
        data[2023]=255;
        data[2022]=255;
        data[2021]=255;
        data[2020]=255;
        data[2019]=255;
        data[2018]=255;
        data[2017]=255;
        data[2016]=255;
        data[2015]=255;
        data[2014]=255;
        data[2013]=255;
        data[2012]=255;
        data[2011]=255;
        data[2010]=255;
        data[2009]=255;
        data[2008]=255;
        data[2007]=255;
        data[2006]=255;
        data[2005]=255;
        data[2004]=255;
        data[2003]=255;
        data[2002]=255;
        data[2001]=255;
        data[2000]=255;
        data[1999]=255;
        data[1998]=255;
        data[1997]=255;
        data[1996]=255;
        data[1995]=255;
        data[1994]=255;
        data[1993]=255;
        data[1992]=255;
        data[1991]=255;
        data[1990]=255;
        data[1989]=255;
        data[1988]=255;
        data[1987]=255;
        data[1986]=255;
        data[1985]=255;
        data[1984]=255;
        data[1983]=255;
        data[1982]=255;
        data[1981]=255;
        data[1980]=255;
        data[1979]=255;
        data[1978]=255;
        data[1977]=255;
        data[1976]=255;
        data[1975]=255;
        data[1974]=255;
        data[1973]=255;
        data[1972]=255;
        data[1971]=255;
        data[1970]=255;
        data[1969]=255;
        data[1968]=255;
        data[1967]=255;
        data[1966]=255;
        data[1965]=255;
        data[1964]=255;
        data[1963]=255;
        data[1962]=255;
        data[1961]=255;
        data[1960]=255;
        data[1959]=255;
        data[1958]=255;
        data[1957]=255;
        data[1956]=255;
        data[1955]=255;
        data[1954]=255;
        data[1953]=255;
        data[1952]=255;
        data[1951]=255;
        data[1950]=255;
        data[1949]=255;
        data[1948]=255;
        data[1947]=255;
        data[1946]=255;
        data[1945]=255;
        data[1944]=255;
        data[1943]=255;
        data[1942]=255;
        data[1941]=255;
        data[1940]=255;
        data[1939]=255;
        data[1938]=255;
        data[1937]=255;
        data[1936]=255;
        data[1935]=255;
        data[1934]=255;
        data[1933]=255;
        data[1932]=255;
        data[1931]=255;
        data[1930]=255;
        data[1929]=255;
        data[1928]=255;
        data[1927]=255;
        data[1926]=255;
        data[1925]=255;
        data[1924]=255;
        data[1923]=255;
        data[1922]=255;
        data[1921]=255;
        data[1920]=255;
        data[1919]=255;
        data[1918]=255;
        data[1917]=255;
        data[1916]=255;
        data[1915]=255;
        data[1914]=255;
        data[1913]=255;
        data[1912]=255;
        data[1911]=255;
        data[1910]=255;
        data[1909]=255;
        data[1908]=255;
        data[1907]=255;
        data[1906]=255;
        data[1905]=255;
        data[1904]=255;
        data[1903]=255;
        data[1902]=255;
        data[1901]=255;
        data[1900]=255;
        data[1899]=255;
        data[1898]=255;
        data[1897]=255;
        data[1896]=255;
        data[1895]=255;
        data[1894]=255;
        data[1893]=255;
        data[1892]=255;
        data[1891]=255;
        data[1890]=255;
        data[1889]=255;
        data[1888]=255;
        data[1887]=255;
        data[1886]=255;
        data[1885]=255;
        data[1884]=255;
        data[1883]=255;
        data[1882]=255;
        data[1881]=255;
        data[1880]=255;
        data[1879]=255;
        data[1878]=255;
        data[1877]=255;
        data[1876]=255;
        data[1875]=255;
        data[1874]=255;
        data[1873]=255;
        data[1872]=255;
        data[1871]=255;
        data[1870]=255;
        data[1869]=255;
        data[1868]=255;
        data[1867]=255;
        data[1866]=255;
        data[1865]=255;
        data[1864]=255;
        data[1863]=255;
        data[1862]=255;
        data[1861]=255;
        data[1860]=255;
        data[1859]=255;
        data[1858]=255;
        data[1857]=255;
        data[1856]=255;
        data[1855]=255;
        data[1854]=255;
        data[1853]=255;
        data[1852]=255;
        data[1851]=255;
        data[1850]=255;
        data[1849]=255;
        data[1848]=255;
        data[1847]=255;
        data[1846]=255;
        data[1845]=255;
        data[1844]=255;
        data[1843]=255;
        data[1842]=255;
        data[1841]=255;
        data[1840]=255;
        data[1839]=255;
        data[1838]=255;
        data[1837]=255;
        data[1836]=255;
        data[1835]=255;
        data[1834]=255;
        data[1833]=255;
        data[1832]=255;
        data[1831]=255;
        data[1830]=255;
        data[1829]=255;
        data[1828]=255;
        data[1827]=255;
        data[1826]=255;
        data[1825]=255;
        data[1824]=255;
        data[1823]=255;
        data[1822]=255;
        data[1821]=255;
        data[1820]=255;
        data[1819]=255;
        data[1818]=255;
        data[1817]=255;
        data[1816]=255;
        data[1815]=255;
        data[1814]=255;
        data[1813]=255;
        data[1812]=255;
        data[1811]=255;
        data[1810]=255;
        data[1809]=255;
        data[1808]=255;
        data[1807]=255;
        data[1806]=255;
        data[1805]=255;
        data[1804]=255;
        data[1803]=255;
        data[1802]=255;
        data[1801]=255;
        data[1800]=255;
        data[1799]=255;
        data[1798]=255;
        data[1797]=255;
        data[1796]=255;
        data[1795]=255;
        data[1794]=255;
        data[1793]=255;
        data[1792]=255;
        data[1791]=255;
        data[1790]=255;
        data[1789]=255;
        data[1788]=255;
        data[1787]=255;
        data[1786]=255;
        data[1785]=255;
        data[1784]=255;
        data[1783]=255;
        data[1782]=255;
        data[1781]=255;
        data[1780]=255;
        data[1779]=255;
        data[1778]=255;
        data[1777]=255;
        data[1776]=255;
        data[1775]=255;
        data[1774]=255;
        data[1773]=255;
        data[1772]=255;
        data[1771]=255;
        data[1770]=255;
        data[1769]=255;
        data[1768]=255;
        data[1767]=255;
        data[1766]=255;
        data[1765]=255;
        data[1764]=255;
        data[1763]=255;
        data[1762]=255;
        data[1761]=255;
        data[1760]=255;
        data[1759]=255;
        data[1758]=255;
        data[1757]=255;
        data[1756]=255;
        data[1755]=255;
        data[1754]=255;
        data[1753]=255;
        data[1752]=255;
        data[1751]=255;
        data[1750]=255;
        data[1749]=255;
        data[1748]=255;
        data[1747]=255;
        data[1746]=255;
        data[1745]=255;
        data[1744]=255;
        data[1743]=255;
        data[1742]=255;
        data[1741]=255;
        data[1740]=255;
        data[1739]=255;
        data[1738]=255;
        data[1737]=255;
        data[1736]=255;
        data[1735]=255;
        data[1734]=255;
        data[1733]=255;
        data[1732]=255;
        data[1731]=255;
        data[1730]=255;
        data[1729]=255;
        data[1728]=255;
        data[1727]=255;
        data[1726]=255;
        data[1725]=255;
        data[1724]=255;
        data[1723]=255;
        data[1722]=255;
        data[1721]=255;
        data[1720]=255;
        data[1719]=255;
        data[1718]=255;
        data[1717]=255;
        data[1716]=255;
        data[1715]=255;
        data[1714]=255;
        data[1713]=255;
        data[1712]=255;
        data[1711]=255;
        data[1710]=255;
        data[1709]=255;
        data[1708]=255;
        data[1707]=255;
        data[1706]=255;
        data[1705]=255;
        data[1704]=255;
        data[1703]=255;
        data[1702]=255;
        data[1701]=255;
        data[1700]=255;
        data[1699]=255;
        data[1698]=255;
        data[1697]=255;
        data[1696]=255;
        data[1695]=255;
        data[1694]=255;
        data[1693]=255;
        data[1692]=255;
        data[1691]=255;
        data[1690]=255;
        data[1689]=255;
        data[1688]=255;
        data[1687]=255;
        data[1686]=255;
        data[1685]=255;
        data[1684]=255;
        data[1683]=255;
        data[1682]=255;
        data[1681]=255;
        data[1680]=255;
        data[1679]=255;
        data[1678]=255;
        data[1677]=255;
        data[1676]=255;
        data[1675]=255;
        data[1674]=255;
        data[1673]=255;
        data[1672]=255;
        data[1671]=255;
        data[1670]=255;
        data[1669]=255;
        data[1668]=255;
        data[1667]=255;
        data[1666]=255;
        data[1665]=255;
        data[1664]=255;
        data[1663]=255;
        data[1662]=255;
        data[1661]=255;
        data[1660]=255;
        data[1659]=255;
        data[1658]=255;
        data[1657]=255;
        data[1656]=255;
        data[1655]=255;
        data[1654]=255;
        data[1653]=255;
        data[1652]=255;
        data[1651]=255;
        data[1650]=255;
        data[1649]=255;
        data[1648]=255;
        data[1647]=255;
        data[1646]=255;
        data[1645]=255;
        data[1644]=255;
        data[1643]=255;
        data[1642]=255;
        data[1641]=255;
        data[1640]=255;
        data[1639]=255;
        data[1638]=255;
        data[1637]=255;
        data[1636]=255;
        data[1635]=255;
        data[1634]=255;
        data[1633]=255;
        data[1632]=255;
        data[1631]=255;
        data[1630]=255;
        data[1629]=255;
        data[1628]=255;
        data[1627]=255;
        data[1626]=255;
        data[1625]=255;
        data[1624]=255;
        data[1623]=255;
        data[1622]=255;
        data[1621]=255;
        data[1620]=255;
        data[1619]=255;
        data[1618]=255;
        data[1617]=255;
        data[1616]=255;
        data[1615]=255;
        data[1614]=255;
        data[1613]=255;
        data[1612]=255;
        data[1611]=255;
        data[1610]=255;
        data[1609]=255;
        data[1608]=255;
        data[1607]=255;
        data[1606]=255;
        data[1605]=255;
        data[1604]=255;
        data[1603]=255;
        data[1602]=255;
        data[1601]=255;
        data[1600]=255;
        data[1599]=255;
        data[1598]=255;
        data[1597]=255;
        data[1596]=255;
        data[1595]=255;
        data[1594]=255;
        data[1593]=255;
        data[1592]=255;
        data[1591]=255;
        data[1590]=255;
        data[1589]=255;
        data[1588]=255;
        data[1587]=255;
        data[1586]=255;
        data[1585]=255;
        data[1584]=255;
        data[1583]=255;
        data[1582]=255;
        data[1581]=255;
        data[1580]=255;
        data[1579]=255;
        data[1578]=255;
        data[1577]=255;
        data[1576]=255;
        data[1575]=255;
        data[1574]=255;
        data[1573]=255;
        data[1572]=255;
        data[1571]=255;
        data[1570]=255;
        data[1569]=255;
        data[1568]=255;
        data[1567]=255;
        data[1566]=255;
        data[1565]=255;
        data[1564]=255;
        data[1563]=255;
        data[1562]=255;
        data[1561]=255;
        data[1560]=255;
        data[1559]=255;
        data[1558]=255;
        data[1557]=255;
        data[1556]=255;
        data[1555]=255;
        data[1554]=255;
        data[1553]=255;
        data[1552]=255;
        data[1551]=255;
        data[1550]=255;
        data[1549]=255;
        data[1548]=255;
        data[1547]=255;
        data[1546]=255;
        data[1545]=255;
        data[1544]=255;
        data[1543]=255;
        data[1542]=255;
        data[1541]=255;
        data[1540]=255;
        data[1539]=255;
        data[1538]=255;
        data[1537]=255;
        data[1536]=255;
        data[1535]=255;
        data[1534]=255;
        data[1533]=255;
        data[1532]=255;
        data[1531]=255;
        data[1530]=255;
        data[1529]=255;
        data[1528]=255;
        data[1527]=255;
        data[1526]=255;
        data[1525]=255;
        data[1524]=255;
        data[1523]=0;
        data[1522]=0;
        data[1521]=0;
        data[1520]=0;
        data[1519]=0;
        data[1518]=0;
        data[1517]=0;
        data[1516]=0;
        data[1515]=0;
        data[1514]=0;
        data[1513]=0;
        data[1512]=0;
        data[1511]=0;
        data[1510]=0;
        data[1509]=0;
        data[1508]=0;
        data[1507]=0;
        data[1506]=0;
        data[1505]=0;
        data[1504]=0;
        data[1503]=0;
        data[1502]=0;
        data[1501]=0;
        data[1500]=0;
        data[1499]=0;
        data[1498]=0;
        data[1497]=0;
        data[1496]=0;
        data[1495]=0;
        data[1494]=0;
        data[1493]=0;
        data[1492]=0;
        data[1491]=0;
        data[1490]=0;
        data[1489]=0;
        data[1488]=0;
        data[1487]=0;
        data[1486]=0;
        data[1485]=0;
        data[1484]=0;
        data[1483]=0;
        data[1482]=0;
        data[1481]=0;
        data[1480]=0;
        data[1479]=0;
        data[1478]=0;
        data[1477]=0;
        data[1476]=0;
        data[1475]=0;
        data[1474]=0;
        data[1473]=0;
        data[1472]=0;
        data[1471]=0;
        data[1470]=0;
        data[1469]=0;
        data[1468]=0;
        data[1467]=0;
        data[1466]=0;
        data[1465]=0;
        data[1464]=0;
        data[1463]=0;
        data[1462]=0;
        data[1461]=0;
        data[1460]=0;
        data[1459]=0;
        data[1458]=0;
        data[1457]=0;
        data[1456]=0;
        data[1455]=0;
        data[1454]=0;
        data[1453]=0;
        data[1452]=0;
        data[1451]=0;
        data[1450]=0;
        data[1449]=0;
        data[1448]=0;
        data[1447]=0;
        data[1446]=0;
        data[1445]=0;
        data[1444]=0;
        data[1443]=0;
        data[1442]=0;
        data[1441]=0;
        data[1440]=0;
        data[1439]=0;
        data[1438]=0;
        data[1437]=0;
        data[1436]=0;
        data[1435]=0;
        data[1434]=0;
        data[1433]=0;
        data[1432]=0;
        data[1431]=0;
        data[1430]=0;
        data[1429]=0;
        data[1428]=0;
        data[1427]=0;
        data[1426]=0;
        data[1425]=0;
        data[1424]=0;
        data[1423]=0;
        data[1422]=0;
        data[1421]=0;
        data[1420]=0;
        data[1419]=0;
        data[1418]=0;
        data[1417]=0;
        data[1416]=0;
        data[1415]=0;
        data[1414]=0;
        data[1413]=0;
        data[1412]=0;
        data[1411]=0;
        data[1410]=0;
        data[1409]=0;
        data[1408]=0;
        data[1407]=0;
        data[1406]=0;
        data[1405]=0;
        data[1404]=0;
        data[1403]=0;
        data[1402]=0;
        data[1401]=0;
        data[1400]=0;
        data[1399]=0;
        data[1398]=0;
        data[1397]=0;
        data[1396]=0;
        data[1395]=0;
        data[1394]=0;
        data[1393]=0;
        data[1392]=0;
        data[1391]=0;
        data[1390]=0;
        data[1389]=0;
        data[1388]=0;
        data[1387]=0;
        data[1386]=0;
        data[1385]=0;
        data[1384]=0;
        data[1383]=0;
        data[1382]=0;
        data[1381]=0;
        data[1380]=0;
        data[1379]=0;
        data[1378]=0;
        data[1377]=0;
        data[1376]=0;
        data[1375]=0;
        data[1374]=0;
        data[1373]=0;
        data[1372]=0;
        data[1371]=0;
        data[1370]=0;
        data[1369]=0;
        data[1368]=0;
        data[1367]=0;
        data[1366]=0;
        data[1365]=0;
        data[1364]=0;
        data[1363]=0;
        data[1362]=0;
        data[1361]=0;
        data[1360]=0;
        data[1359]=0;
        data[1358]=0;
        data[1357]=0;
        data[1356]=0;
        data[1355]=0;
        data[1354]=0;
        data[1353]=0;
        data[1352]=0;
        data[1351]=0;
        data[1350]=0;
        data[1349]=0;
        data[1348]=0;
        data[1347]=0;
        data[1346]=0;
        data[1345]=0;
        data[1344]=0;
        data[1343]=0;
        data[1342]=0;
        data[1341]=0;
        data[1340]=0;
        data[1339]=0;
        data[1338]=0;
        data[1337]=0;
        data[1336]=0;
        data[1335]=0;
        data[1334]=0;
        data[1333]=0;
        data[1332]=0;
        data[1331]=0;
        data[1330]=0;
        data[1329]=0;
        data[1328]=0;
        data[1327]=0;
        data[1326]=0;
        data[1325]=0;
        data[1324]=0;
        data[1323]=0;
        data[1322]=0;
        data[1321]=0;
        data[1320]=0;
        data[1319]=0;
        data[1318]=0;
        data[1317]=0;
        data[1316]=0;
        data[1315]=0;
        data[1314]=0;
        data[1313]=0;
        data[1312]=0;
        data[1311]=0;
        data[1310]=0;
        data[1309]=0;
        data[1308]=0;
        data[1307]=0;
        data[1306]=0;
        data[1305]=0;
        data[1304]=0;
        data[1303]=0;
        data[1302]=0;
        data[1301]=0;
        data[1300]=0;
        data[1299]=0;
        data[1298]=0;
        data[1297]=0;
        data[1296]=0;
        data[1295]=0;
        data[1294]=0;
        data[1293]=0;
        data[1292]=0;
        data[1291]=0;
        data[1290]=0;
        data[1289]=0;
        data[1288]=0;
        data[1287]=0;
        data[1286]=0;
        data[1285]=0;
        data[1284]=0;
        data[1283]=0;
        data[1282]=0;
        data[1281]=0;
        data[1280]=0;
        data[1279]=0;
        data[1278]=0;
        data[1277]=0;
        data[1276]=0;
        data[1275]=0;
        data[1274]=0;
        data[1273]=0;
        data[1272]=0;
        data[1271]=0;
        data[1270]=0;
        data[1269]=0;
        data[1268]=0;
        data[1267]=0;
        data[1266]=0;
        data[1265]=0;
        data[1264]=0;
        data[1263]=0;
        data[1262]=0;
        data[1261]=0;
        data[1260]=0;
        data[1259]=0;
        data[1258]=0;
        data[1257]=0;
        data[1256]=0;
        data[1255]=0;
        data[1254]=0;
        data[1253]=0;
        data[1252]=0;
        data[1251]=0;
        data[1250]=0;
        data[1249]=0;
        data[1248]=0;
        data[1247]=0;
        data[1246]=0;
        data[1245]=0;
        data[1244]=0;
        data[1243]=0;
        data[1242]=0;
        data[1241]=0;
        data[1240]=0;
        data[1239]=0;
        data[1238]=0;
        data[1237]=0;
        data[1236]=0;
        data[1235]=0;
        data[1234]=0;
        data[1233]=0;
        data[1232]=0;
        data[1231]=0;
        data[1230]=0;
        data[1229]=0;
        data[1228]=0;
        data[1227]=0;
        data[1226]=0;
        data[1225]=0;
        data[1224]=0;
        data[1223]=0;
        data[1222]=0;
        data[1221]=0;
        data[1220]=0;
        data[1219]=0;
        data[1218]=0;
        data[1217]=0;
        data[1216]=0;
        data[1215]=0;
        data[1214]=0;
        data[1213]=0;
        data[1212]=0;
        data[1211]=0;
        data[1210]=0;
        data[1209]=0;
        data[1208]=0;
        data[1207]=0;
        data[1206]=0;
        data[1205]=0;
        data[1204]=0;
        data[1203]=0;
        data[1202]=0;
        data[1201]=0;
        data[1200]=0;
        data[1199]=0;
        data[1198]=0;
        data[1197]=0;
        data[1196]=0;
        data[1195]=0;
        data[1194]=0;
        data[1193]=0;
        data[1192]=0;
        data[1191]=0;
        data[1190]=0;
        data[1189]=0;
        data[1188]=0;
        data[1187]=0;
        data[1186]=0;
        data[1185]=0;
        data[1184]=0;
        data[1183]=0;
        data[1182]=0;
        data[1181]=0;
        data[1180]=0;
        data[1179]=0;
        data[1178]=0;
        data[1177]=0;
        data[1176]=0;
        data[1175]=0;
        data[1174]=0;
        data[1173]=0;
        data[1172]=0;
        data[1171]=0;
        data[1170]=0;
        data[1169]=0;
        data[1168]=0;
        data[1167]=0;
        data[1166]=0;
        data[1165]=0;
        data[1164]=0;
        data[1163]=0;
        data[1162]=0;
        data[1161]=0;
        data[1160]=0;
        data[1159]=0;
        data[1158]=0;
        data[1157]=0;
        data[1156]=0;
        data[1155]=0;
        data[1154]=0;
        data[1153]=0;
        data[1152]=0;
        data[1151]=0;
        data[1150]=0;
        data[1149]=0;
        data[1148]=0;
        data[1147]=0;
        data[1146]=0;
        data[1145]=0;
        data[1144]=0;
        data[1143]=0;
        data[1142]=0;
        data[1141]=0;
        data[1140]=0;
        data[1139]=0;
        data[1138]=0;
        data[1137]=0;
        data[1136]=0;
        data[1135]=0;
        data[1134]=0;
        data[1133]=0;
        data[1132]=0;
        data[1131]=0;
        data[1130]=0;
        data[1129]=0;
        data[1128]=0;
        data[1127]=0;
        data[1126]=0;
        data[1125]=0;
        data[1124]=0;
        data[1123]=0;
        data[1122]=0;
        data[1121]=0;
        data[1120]=0;
        data[1119]=0;
        data[1118]=0;
        data[1117]=0;
        data[1116]=0;
        data[1115]=0;
        data[1114]=0;
        data[1113]=0;
        data[1112]=0;
        data[1111]=0;
        data[1110]=0;
        data[1109]=0;
        data[1108]=0;
        data[1107]=0;
        data[1106]=0;
        data[1105]=0;
        data[1104]=0;
        data[1103]=0;
        data[1102]=0;
        data[1101]=0;
        data[1100]=0;
        data[1099]=0;
        data[1098]=0;
        data[1097]=0;
        data[1096]=0;
        data[1095]=0;
        data[1094]=0;
        data[1093]=0;
        data[1092]=0;
        data[1091]=0;
        data[1090]=0;
        data[1089]=0;
        data[1088]=0;
        data[1087]=0;
        data[1086]=0;
        data[1085]=0;
        data[1084]=0;
        data[1083]=0;
        data[1082]=0;
        data[1081]=0;
        data[1080]=0;
        data[1079]=0;
        data[1078]=0;
        data[1077]=0;
        data[1076]=0;
        data[1075]=0;
        data[1074]=0;
        data[1073]=0;
        data[1072]=0;
        data[1071]=0;
        data[1070]=0;
        data[1069]=0;
        data[1068]=0;
        data[1067]=0;
        data[1066]=0;
        data[1065]=0;
        data[1064]=0;
        data[1063]=0;
        data[1062]=0;
        data[1061]=0;
        data[1060]=0;
        data[1059]=0;
        data[1058]=0;
        data[1057]=0;
        data[1056]=0;
        data[1055]=0;
        data[1054]=0;
        data[1053]=0;
        data[1052]=0;
        data[1051]=0;
        data[1050]=0;
        data[1049]=0;
        data[1048]=0;
        data[1047]=0;
        data[1046]=0;
        data[1045]=0;
        data[1044]=0;
        data[1043]=0;
        data[1042]=0;
        data[1041]=0;
        data[1040]=0;
        data[1039]=0;
        data[1038]=0;
        data[1037]=0;
        data[1036]=0;
        data[1035]=0;
        data[1034]=0;
        data[1033]=0;
        data[1032]=0;
        data[1031]=0;
        data[1030]=0;
        data[1029]=0;
        data[1028]=0;
        data[1027]=0;
        data[1026]=0;
        data[1025]=0;
        data[1024]=0;
        data[1023]=0;
        data[1022]=0;
        data[1021]=0;
        data[1020]=0;
        data[1019]=0;
        data[1018]=0;
        data[1017]=0;
        data[1016]=0;
        data[1015]=0;
        data[1014]=0;
        data[1013]=0;
        data[1012]=0;
        data[1011]=0;
        data[1010]=0;
        data[1009]=0;
        data[1008]=0;
        data[1007]=0;
        data[1006]=0;
        data[1005]=0;
        data[1004]=0;
        data[1003]=0;
        data[1002]=0;
        data[1001]=0;
        data[1000]=0;
        data[999]=126;
        data[998]=125;
        data[997]=125;
        data[996]=124;
        data[995]=123;
        data[994]=122;
        data[993]=121;
        data[992]=121;
        data[991]=120;
        data[990]=119;
        data[989]=118;
        data[988]=117;
        data[987]=117;
        data[986]=116;
        data[985]=115;
        data[984]=114;
        data[983]=113;
        data[982]=113;
        data[981]=112;
        data[980]=111;
        data[979]=110;
        data[978]=109;
        data[977]=109;
        data[976]=108;
        data[975]=107;
        data[974]=106;
        data[973]=105;
        data[972]=105;
        data[971]=104;
        data[970]=103;
        data[969]=102;
        data[968]=101;
        data[967]=101;
        data[966]=100;
        data[965]=99;
        data[964]=98;
        data[963]=98;
        data[962]=97;
        data[961]=96;
        data[960]=95;
        data[959]=94;
        data[958]=94;
        data[957]=93;
        data[956]=92;
        data[955]=91;
        data[954]=91;
        data[953]=90;
        data[952]=89;
        data[951]=88;
        data[950]=87;
        data[949]=87;
        data[948]=86;
        data[947]=85;
        data[946]=84;
        data[945]=84;
        data[944]=83;
        data[943]=82;
        data[942]=81;
        data[941]=81;
        data[940]=80;
        data[939]=79;
        data[938]=78;
        data[937]=78;
        data[936]=77;
        data[935]=76;
        data[934]=75;
        data[933]=75;
        data[932]=74;
        data[931]=73;
        data[930]=73;
        data[929]=72;
        data[928]=71;
        data[927]=70;
        data[926]=70;
        data[925]=69;
        data[924]=68;
        data[923]=67;
        data[922]=67;
        data[921]=66;
        data[920]=65;
        data[919]=65;
        data[918]=64;
        data[917]=63;
        data[916]=63;
        data[915]=62;
        data[914]=61;
        data[913]=60;
        data[912]=60;
        data[911]=59;
        data[910]=58;
        data[909]=58;
        data[908]=57;
        data[907]=56;
        data[906]=56;
        data[905]=55;
        data[904]=54;
        data[903]=54;
        data[902]=53;
        data[901]=52;
        data[900]=52;
        data[899]=51;
        data[898]=50;
        data[897]=50;
        data[896]=49;
        data[895]=49;
        data[894]=48;
        data[893]=47;
        data[892]=47;
        data[891]=46;
        data[890]=45;
        data[889]=45;
        data[888]=44;
        data[887]=44;
        data[886]=43;
        data[885]=42;
        data[884]=42;
        data[883]=41;
        data[882]=41;
        data[881]=40;
        data[880]=39;
        data[879]=39;
        data[878]=38;
        data[877]=38;
        data[876]=37;
        data[875]=36;
        data[874]=36;
        data[873]=35;
        data[872]=35;
        data[871]=34;
        data[870]=34;
        data[869]=33;
        data[868]=33;
        data[867]=32;
        data[866]=32;
        data[865]=31;
        data[864]=30;
        data[863]=30;
        data[862]=29;
        data[861]=29;
        data[860]=28;
        data[859]=28;
        data[858]=27;
        data[857]=27;
        data[856]=26;
        data[855]=26;
        data[854]=25;
        data[853]=25;
        data[852]=24;
        data[851]=24;
        data[850]=23;
        data[849]=23;
        data[848]=23;
        data[847]=22;
        data[846]=22;
        data[845]=21;
        data[844]=21;
        data[843]=20;
        data[842]=20;
        data[841]=19;
        data[840]=19;
        data[839]=18;
        data[838]=18;
        data[837]=18;
        data[836]=17;
        data[835]=17;
        data[834]=16;
        data[833]=16;
        data[832]=16;
        data[831]=15;
        data[830]=15;
        data[829]=14;
        data[828]=14;
        data[827]=14;
        data[826]=13;
        data[825]=13;
        data[824]=13;
        data[823]=12;
        data[822]=12;
        data[821]=12;
        data[820]=11;
        data[819]=11;
        data[818]=11;
        data[817]=10;
        data[816]=10;
        data[815]=10;
        data[814]=9;
        data[813]=9;
        data[812]=9;
        data[811]=8;
        data[810]=8;
        data[809]=8;
        data[808]=7;
        data[807]=7;
        data[806]=7;
        data[805]=7;
        data[804]=6;
        data[803]=6;
        data[802]=6;
        data[801]=6;
        data[800]=5;
        data[799]=5;
        data[798]=5;
        data[797]=5;
        data[796]=4;
        data[795]=4;
        data[794]=4;
        data[793]=4;
        data[792]=3;
        data[791]=3;
        data[790]=3;
        data[789]=3;
        data[788]=3;
        data[787]=2;
        data[786]=2;
        data[785]=2;
        data[784]=2;
        data[783]=2;
        data[782]=2;
        data[781]=1;
        data[780]=1;
        data[779]=1;
        data[778]=1;
        data[777]=1;
        data[776]=1;
        data[775]=1;
        data[774]=0;
        data[773]=0;
        data[772]=0;
        data[771]=0;
        data[770]=0;
        data[769]=0;
        data[768]=0;
        data[767]=0;
        data[766]=0;
        data[765]=0;
        data[764]=0;
        data[763]=0;
        data[762]=0;
        data[761]=0;
        data[760]=0;
        data[759]=0;
        data[758]=0;
        data[757]=0;
        data[756]=0;
        data[755]=0;
        data[754]=0;
        data[753]=0;
        data[752]=0;
        data[751]=0;
        data[750]=0;
        data[749]=0;
        data[748]=0;
        data[747]=0;
        data[746]=0;
        data[745]=0;
        data[744]=0;
        data[743]=0;
        data[742]=0;
        data[741]=0;
        data[740]=0;
        data[739]=0;
        data[738]=0;
        data[737]=0;
        data[736]=0;
        data[735]=0;
        data[734]=0;
        data[733]=0;
        data[732]=0;
        data[731]=0;
        data[730]=0;
        data[729]=0;
        data[728]=0;
        data[727]=0;
        data[726]=0;
        data[725]=1;
        data[724]=1;
        data[723]=1;
        data[722]=1;
        data[721]=1;
        data[720]=1;
        data[719]=1;
        data[718]=2;
        data[717]=2;
        data[716]=2;
        data[715]=2;
        data[714]=2;
        data[713]=2;
        data[712]=3;
        data[711]=3;
        data[710]=3;
        data[709]=3;
        data[708]=3;
        data[707]=4;
        data[706]=4;
        data[705]=4;
        data[704]=4;
        data[703]=5;
        data[702]=5;
        data[701]=5;
        data[700]=5;
        data[699]=6;
        data[698]=6;
        data[697]=6;
        data[696]=6;
        data[695]=7;
        data[694]=7;
        data[693]=7;
        data[692]=7;
        data[691]=8;
        data[690]=8;
        data[689]=8;
        data[688]=9;
        data[687]=9;
        data[686]=9;
        data[685]=10;
        data[684]=10;
        data[683]=10;
        data[682]=11;
        data[681]=11;
        data[680]=11;
        data[679]=12;
        data[678]=12;
        data[677]=12;
        data[676]=13;
        data[675]=13;
        data[674]=13;
        data[673]=14;
        data[672]=14;
        data[671]=14;
        data[670]=15;
        data[669]=15;
        data[668]=16;
        data[667]=16;
        data[666]=16;
        data[665]=17;
        data[664]=17;
        data[663]=18;
        data[662]=18;
        data[661]=18;
        data[660]=19;
        data[659]=19;
        data[658]=20;
        data[657]=20;
        data[656]=21;
        data[655]=21;
        data[654]=22;
        data[653]=22;
        data[652]=23;
        data[651]=23;
        data[650]=23;
        data[649]=24;
        data[648]=24;
        data[647]=25;
        data[646]=25;
        data[645]=26;
        data[644]=26;
        data[643]=27;
        data[642]=27;
        data[641]=28;
        data[640]=28;
        data[639]=29;
        data[638]=29;
        data[637]=30;
        data[636]=30;
        data[635]=31;
        data[634]=32;
        data[633]=32;
        data[632]=33;
        data[631]=33;
        data[630]=34;
        data[629]=34;
        data[628]=35;
        data[627]=35;
        data[626]=36;
        data[625]=36;
        data[624]=37;
        data[623]=38;
        data[622]=38;
        data[621]=39;
        data[620]=39;
        data[619]=40;
        data[618]=41;
        data[617]=41;
        data[616]=42;
        data[615]=42;
        data[614]=43;
        data[613]=44;
        data[612]=44;
        data[611]=45;
        data[610]=45;
        data[609]=46;
        data[608]=47;
        data[607]=47;
        data[606]=48;
        data[605]=49;
        data[604]=49;
        data[603]=50;
        data[602]=50;
        data[601]=51;
        data[600]=52;
        data[599]=52;
        data[598]=53;
        data[597]=54;
        data[596]=54;
        data[595]=55;
        data[594]=56;
        data[593]=56;
        data[592]=57;
        data[591]=58;
        data[590]=58;
        data[589]=59;
        data[588]=60;
        data[587]=60;
        data[586]=61;
        data[585]=62;
        data[584]=63;
        data[583]=63;
        data[582]=64;
        data[581]=65;
        data[580]=65;
        data[579]=66;
        data[578]=67;
        data[577]=67;
        data[576]=68;
        data[575]=69;
        data[574]=70;
        data[573]=70;
        data[572]=71;
        data[571]=72;
        data[570]=73;
        data[569]=73;
        data[568]=74;
        data[567]=75;
        data[566]=75;
        data[565]=76;
        data[564]=77;
        data[563]=78;
        data[562]=78;
        data[561]=79;
        data[560]=80;
        data[559]=81;
        data[558]=81;
        data[557]=82;
        data[556]=83;
        data[555]=84;
        data[554]=84;
        data[553]=85;
        data[552]=86;
        data[551]=87;
        data[550]=87;
        data[549]=88;
        data[548]=89;
        data[547]=90;
        data[546]=91;
        data[545]=91;
        data[544]=92;
        data[543]=93;
        data[542]=94;
        data[541]=94;
        data[540]=95;
        data[539]=96;
        data[538]=97;
        data[537]=98;
        data[536]=98;
        data[535]=99;
        data[534]=100;
        data[533]=101;
        data[532]=101;
        data[531]=102;
        data[530]=103;
        data[529]=104;
        data[528]=105;
        data[527]=105;
        data[526]=106;
        data[525]=107;
        data[524]=108;
        data[523]=109;
        data[522]=109;
        data[521]=110;
        data[520]=111;
        data[519]=112;
        data[518]=113;
        data[517]=113;
        data[516]=114;
        data[515]=115;
        data[514]=116;
        data[513]=117;
        data[512]=117;
        data[511]=118;
        data[510]=119;
        data[509]=120;
        data[508]=121;
        data[507]=121;
        data[506]=122;
        data[505]=123;
        data[504]=124;
        data[503]=125;
        data[502]=125;
        data[501]=126;
        data[500]=127;
        data[499]=128;
        data[498]=129;
        data[497]=129;
        data[496]=130;
        data[495]=131;
        data[494]=132;
        data[493]=133;
        data[492]=133;
        data[491]=134;
        data[490]=135;
        data[489]=136;
        data[488]=137;
        data[487]=137;
        data[486]=138;
        data[485]=139;
        data[484]=140;
        data[483]=141;
        data[482]=141;
        data[481]=142;
        data[480]=143;
        data[479]=144;
        data[478]=145;
        data[477]=145;
        data[476]=146;
        data[475]=147;
        data[474]=148;
        data[473]=149;
        data[472]=149;
        data[471]=150;
        data[470]=151;
        data[469]=152;
        data[468]=153;
        data[467]=153;
        data[466]=154;
        data[465]=155;
        data[464]=156;
        data[463]=156;
        data[462]=157;
        data[461]=158;
        data[460]=159;
        data[459]=160;
        data[458]=160;
        data[457]=161;
        data[456]=162;
        data[455]=163;
        data[454]=163;
        data[453]=164;
        data[452]=165;
        data[451]=166;
        data[450]=167;
        data[449]=167;
        data[448]=168;
        data[447]=169;
        data[446]=170;
        data[445]=170;
        data[444]=171;
        data[443]=172;
        data[442]=173;
        data[441]=173;
        data[440]=174;
        data[439]=175;
        data[438]=176;
        data[437]=176;
        data[436]=177;
        data[435]=178;
        data[434]=179;
        data[433]=179;
        data[432]=180;
        data[431]=181;
        data[430]=181;
        data[429]=182;
        data[428]=183;
        data[427]=184;
        data[426]=184;
        data[425]=185;
        data[424]=186;
        data[423]=187;
        data[422]=187;
        data[421]=188;
        data[420]=189;
        data[419]=189;
        data[418]=190;
        data[417]=191;
        data[416]=191;
        data[415]=192;
        data[414]=193;
        data[413]=194;
        data[412]=194;
        data[411]=195;
        data[410]=196;
        data[409]=196;
        data[408]=197;
        data[407]=198;
        data[406]=198;
        data[405]=199;
        data[404]=200;
        data[403]=200;
        data[402]=201;
        data[401]=202;
        data[400]=202;
        data[399]=203;
        data[398]=204;
        data[397]=204;
        data[396]=205;
        data[395]=205;
        data[394]=206;
        data[393]=207;
        data[392]=207;
        data[391]=208;
        data[390]=209;
        data[389]=209;
        data[388]=210;
        data[387]=210;
        data[386]=211;
        data[385]=212;
        data[384]=212;
        data[383]=213;
        data[382]=213;
        data[381]=214;
        data[380]=215;
        data[379]=215;
        data[378]=216;
        data[377]=216;
        data[376]=217;
        data[375]=218;
        data[374]=218;
        data[373]=219;
        data[372]=219;
        data[371]=220;
        data[370]=220;
        data[369]=221;
        data[368]=221;
        data[367]=222;
        data[366]=222;
        data[365]=223;
        data[364]=224;
        data[363]=224;
        data[362]=225;
        data[361]=225;
        data[360]=226;
        data[359]=226;
        data[358]=227;
        data[357]=227;
        data[356]=228;
        data[355]=228;
        data[354]=229;
        data[353]=229;
        data[352]=230;
        data[351]=230;
        data[350]=231;
        data[349]=231;
        data[348]=231;
        data[347]=232;
        data[346]=232;
        data[345]=233;
        data[344]=233;
        data[343]=234;
        data[342]=234;
        data[341]=235;
        data[340]=235;
        data[339]=236;
        data[338]=236;
        data[337]=236;
        data[336]=237;
        data[335]=237;
        data[334]=238;
        data[333]=238;
        data[332]=238;
        data[331]=239;
        data[330]=239;
        data[329]=240;
        data[328]=240;
        data[327]=240;
        data[326]=241;
        data[325]=241;
        data[324]=241;
        data[323]=242;
        data[322]=242;
        data[321]=242;
        data[320]=243;
        data[319]=243;
        data[318]=243;
        data[317]=244;
        data[316]=244;
        data[315]=244;
        data[314]=245;
        data[313]=245;
        data[312]=245;
        data[311]=246;
        data[310]=246;
        data[309]=246;
        data[308]=247;
        data[307]=247;
        data[306]=247;
        data[305]=247;
        data[304]=248;
        data[303]=248;
        data[302]=248;
        data[301]=248;
        data[300]=249;
        data[299]=249;
        data[298]=249;
        data[297]=249;
        data[296]=250;
        data[295]=250;
        data[294]=250;
        data[293]=250;
        data[292]=251;
        data[291]=251;
        data[290]=251;
        data[289]=251;
        data[288]=251;
        data[287]=252;
        data[286]=252;
        data[285]=252;
        data[284]=252;
        data[283]=252;
        data[282]=252;
        data[281]=253;
        data[280]=253;
        data[279]=253;
        data[278]=253;
        data[277]=253;
        data[276]=253;
        data[275]=253;
        data[274]=254;
        data[273]=254;
        data[272]=254;
        data[271]=254;
        data[270]=254;
        data[269]=254;
        data[268]=254;
        data[267]=254;
        data[266]=254;
        data[265]=254;
        data[264]=255;
        data[263]=255;
        data[262]=255;
        data[261]=255;
        data[260]=255;
        data[259]=255;
        data[258]=255;
        data[257]=255;
        data[256]=255;
        data[255]=255;
        data[254]=255;
        data[253]=255;
        data[252]=255;
        data[251]=255;
        data[250]=255;
        data[249]=255;
        data[248]=255;
        data[247]=255;
        data[246]=255;
        data[245]=255;
        data[244]=255;
        data[243]=255;
        data[242]=255;
        data[241]=255;
        data[240]=255;
        data[239]=255;
        data[238]=255;
        data[237]=255;
        data[236]=255;
        data[235]=254;
        data[234]=254;
        data[233]=254;
        data[232]=254;
        data[231]=254;
        data[230]=254;
        data[229]=254;
        data[228]=254;
        data[227]=254;
        data[226]=254;
        data[225]=253;
        data[224]=253;
        data[223]=253;
        data[222]=253;
        data[221]=253;
        data[220]=253;
        data[219]=253;
        data[218]=252;
        data[217]=252;
        data[216]=252;
        data[215]=252;
        data[214]=252;
        data[213]=252;
        data[212]=251;
        data[211]=251;
        data[210]=251;
        data[209]=251;
        data[208]=251;
        data[207]=250;
        data[206]=250;
        data[205]=250;
        data[204]=250;
        data[203]=249;
        data[202]=249;
        data[201]=249;
        data[200]=249;
        data[199]=248;
        data[198]=248;
        data[197]=248;
        data[196]=248;
        data[195]=247;
        data[194]=247;
        data[193]=247;
        data[192]=247;
        data[191]=246;
        data[190]=246;
        data[189]=246;
        data[188]=245;
        data[187]=245;
        data[186]=245;
        data[185]=244;
        data[184]=244;
        data[183]=244;
        data[182]=243;
        data[181]=243;
        data[180]=243;
        data[179]=242;
        data[178]=242;
        data[177]=242;
        data[176]=241;
        data[175]=241;
        data[174]=241;
        data[173]=240;
        data[172]=240;
        data[171]=240;
        data[170]=239;
        data[169]=239;
        data[168]=238;
        data[167]=238;
        data[166]=238;
        data[165]=237;
        data[164]=237;
        data[163]=236;
        data[162]=236;
        data[161]=236;
        data[160]=235;
        data[159]=235;
        data[158]=234;
        data[157]=234;
        data[156]=233;
        data[155]=233;
        data[154]=232;
        data[153]=232;
        data[152]=231;
        data[151]=231;
        data[150]=231;
        data[149]=230;
        data[148]=230;
        data[147]=229;
        data[146]=229;
        data[145]=228;
        data[144]=228;
        data[143]=227;
        data[142]=227;
        data[141]=226;
        data[140]=226;
        data[139]=225;
        data[138]=225;
        data[137]=224;
        data[136]=224;
        data[135]=223;
        data[134]=222;
        data[133]=222;
        data[132]=221;
        data[131]=221;
        data[130]=220;
        data[129]=220;
        data[128]=219;
        data[127]=219;
        data[126]=218;
        data[125]=218;
        data[124]=217;
        data[123]=216;
        data[122]=216;
        data[121]=215;
        data[120]=215;
        data[119]=214;
        data[118]=213;
        data[117]=213;
        data[116]=212;
        data[115]=212;
        data[114]=211;
        data[113]=210;
        data[112]=210;
        data[111]=209;
        data[110]=209;
        data[109]=208;
        data[108]=207;
        data[107]=207;
        data[106]=206;
        data[105]=205;
        data[104]=205;
        data[103]=204;
        data[102]=204;
        data[101]=203;
        data[100]=202;
        data[99]=202;
        data[98]=201;
        data[97]=200;
        data[96]=200;
        data[95]=199;
        data[94]=198;
        data[93]=198;
        data[92]=197;
        data[91]=196;
        data[90]=196;
        data[89]=195;
        data[88]=194;
        data[87]=194;
        data[86]=193;
        data[85]=192;
        data[84]=191;
        data[83]=191;
        data[82]=190;
        data[81]=189;
        data[80]=189;
        data[79]=188;
        data[78]=187;
        data[77]=187;
        data[76]=186;
        data[75]=185;
        data[74]=184;
        data[73]=184;
        data[72]=183;
        data[71]=182;
        data[70]=181;
        data[69]=181;
        data[68]=180;
        data[67]=179;
        data[66]=179;
        data[65]=178;
        data[64]=177;
        data[63]=176;
        data[62]=176;
        data[61]=175;
        data[60]=174;
        data[59]=173;
        data[58]=173;
        data[57]=172;
        data[56]=171;
        data[55]=170;
        data[54]=170;
        data[53]=169;
        data[52]=168;
        data[51]=167;
        data[50]=167;
        data[49]=166;
        data[48]=165;
        data[47]=164;
        data[46]=163;
        data[45]=163;
        data[44]=162;
        data[43]=161;
        data[42]=160;
        data[41]=160;
        data[40]=159;
        data[39]=158;
        data[38]=157;
        data[37]=156;
        data[36]=156;
        data[35]=155;
        data[34]=154;
        data[33]=153;
        data[32]=153;
        data[31]=152;
        data[30]=151;
        data[29]=150;
        data[28]=149;
        data[27]=149;
        data[26]=148;
        data[25]=147;
        data[24]=146;
        data[23]=145;
        data[22]=145;
        data[21]=144;
        data[20]=143;
        data[19]=142;
        data[18]=141;
        data[17]=141;
        data[16]=140;
        data[15]=139;
        data[14]=138;
        data[13]=137;
        data[12]=137;
        data[11]=136;
        data[10]=135;
        data[9]=134;
        data[8]=133;
        data[7]=133;
        data[6]=132;
        data[5]=131;
        data[4]=130;
        data[3]=129;
        data[2]=129;
        data[1]=128;
        data[0]=127;

    end
    always @(posedge clk) begin
        
         otp<=data[{choose,count}];
        count<=(count+1'b1)%mod;
    end
    always @(posedge clk) begin
        if(count==999) cout<=1;
        else cout<=0;
    end
endmodule